--  network.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity network is
		generic(
			N : natural := 321;
			N_SIGNALS : natural := 79;
			N_ROUTES : natural := 91;
			N_LEVELCROSSINGS : natural := 2;
			N_SINGLESWITCHES : natural := 21;
			N_DOUBLEWITCHES : natural := 1;
			N_TRACKCIRCUITS : natural := 47
		);
		port(
			clock : in std_logic;
			processing : in std_logic;
			processed : out std_logic;
			ocupation : in std_logic_vector(N_TRACKCIRCUITS-1 downto 0);
			signals_i : in signals_type;
			signals_o : out signals_type;
			routes_i : in std_logic_vector(N_ROUTES-1 downto 0);
			routes_o : out std_logic_vector(N_ROUTES-1 downto 0);
			levelCrossings_i : in std_logic_vector(N_LEVELCROSSINGS-1 downto 0);
			levelCrossings_o : out std_logic_vector(N_LEVELCROSSINGS-1 downto 0);
			singleSwitches_i : in std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			singleSwitches_o : out std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			doubleSwitches_i : in dSwitches_type;
			doubleSwitches_o : out dSwitches_type;
			reset : in std_logic
		);
	end entity network;
architecture Behavioral of network is
	component levelCrossing_0 is
		port(
			clock : in std_logic;
			ocupation_ne98 : in std_logic;
			ocupation_ne996 : in std_logic;
			ocupation_ne99 : in std_logic;
			R30_command : in routeCommands;
			R31_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc01 : out levelCrossingStates
		);
	end component levelCrossing_0;
	component levelCrossing_1 is
		port(
			clock : in std_logic;
			ocupation_ne98 : in std_logic;
			ocupation_ne996 : in std_logic;
			ocupation_ne99 : in std_logic;
			R30_command : in routeCommands;
			R31_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc02 : out levelCrossingStates
		);
	end component levelCrossing_1;
	component levelCrossing_2 is
		port(
			clock : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne992 : in std_logic;
			ocupation_ne101 : in std_logic;
			R32_command : in routeCommands;
			R33_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc03 : out levelCrossingStates
		);
	end component levelCrossing_2;
	component levelCrossing_3 is
		port(
			clock : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne992 : in std_logic;
			ocupation_ne101 : in std_logic;
			R32_command : in routeCommands;
			R34_command : in routeCommands;
			R35_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc04 : out levelCrossingStates
		);
	end component levelCrossing_3;
	component levelCrossing_4 is
		port(
			clock : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne992 : in std_logic;
			ocupation_ne101 : in std_logic;
			R32_command : in routeCommands;
			R33_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc05 : out levelCrossingStates
		);
	end component levelCrossing_4;
	component levelCrossing_5 is
		port(
			clock : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne992 : in std_logic;
			ocupation_ne101 : in std_logic;
			R32_command : in routeCommands;
			R34_command : in routeCommands;
			R35_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc06 : out levelCrossingStates
		);
	end component levelCrossing_5;
	component singleSwitch_0 is
		port(
			clock : in std_logic;
			R20_command : in routeCommands;
			R41_command : in routeCommands;
			R42_command : in routeCommands;
			R43_command : in routeCommands;
			R49_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D01 : out singleSwitchStates
		);
	end component singleSwitch_0;
	component singleSwitch_1 is
		port(
			clock : in std_logic;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			R58_command : in routeCommands;
			R69_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D08 : out singleSwitchStates
		);
	end component singleSwitch_1;
	component singleSwitch_2 is
		port(
			clock : in std_logic;
			R36_command : in routeCommands;
			R37_command : in routeCommands;
			R38_command : in routeCommands;
			R55_command : in routeCommands;
			R69_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D05 : out singleSwitchStates
		);
	end component singleSwitch_2;
	component singleSwitch_3 is
		port(
			clock : in std_logic;
			R4_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D18 : out singleSwitchStates
		);
	end component singleSwitch_3;
	component singleSwitch_4 is
		port(
			clock : in std_logic;
			R65_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw01 : out singleSwitchStates
		);
	end component singleSwitch_4;
	component singleSwitch_5 is
		port(
			clock : in std_logic;
			R59_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			R82_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D10 : out singleSwitchStates
		);
	end component singleSwitch_5;
	component singleSwitch_6 is
		port(
			clock : in std_logic;
			R26_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			R59_command : in routeCommands;
			R82_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D09 : out singleSwitchStates
		);
	end component singleSwitch_6;
	component singleSwitch_7 is
		port(
			clock : in std_logic;
			R8_command : in routeCommands;
			R28_command : in routeCommands;
			R80_command : in routeCommands;
			R81_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D20 : out singleSwitchStates
		);
	end component singleSwitch_7;
	component singleSwitch_8 is
		port(
			clock : in std_logic;
			R27_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			R78_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D23 : out singleSwitchStates
		);
	end component singleSwitch_8;
	component singleSwitch_9 is
		port(
			clock : in std_logic;
			R43_command : in routeCommands;
			R45_command : in routeCommands;
			R46_command : in routeCommands;
			R49_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D03 : out singleSwitchStates
		);
	end component singleSwitch_9;
	component singleSwitch_10 is
		port(
			clock : in std_logic;
			R2_command : in routeCommands;
			R22_command : in routeCommands;
			R66_command : in routeCommands;
			R67_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D14 : out singleSwitchStates
		);
	end component singleSwitch_10;
	component singleSwitch_11 is
		port(
			clock : in std_logic;
			R21_command : in routeCommands;
			R89_command : in routeCommands;
			R90_command : in routeCommands;
			R91_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw04 : out singleSwitchStates
		);
	end component singleSwitch_11;
	component singleSwitch_12 is
		port(
			clock : in std_logic;
			R11_command : in routeCommands;
			R44_command : in routeCommands;
			R47_command : in routeCommands;
			R50_command : in routeCommands;
			R51_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D04 : out singleSwitchStates
		);
	end component singleSwitch_12;
	component singleSwitch_13 is
		port(
			clock : in std_logic;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			R89_command : in routeCommands;
			R91_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw03 : out singleSwitchStates
		);
	end component singleSwitch_13;
	component singleSwitch_14 is
		port(
			clock : in std_logic;
			R2_command : in routeCommands;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			R67_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D15 : out singleSwitchStates
		);
	end component singleSwitch_14;
	component singleSwitch_15 is
		port(
			clock : in std_logic;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			R65_command : in routeCommands;
			R86_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw02 : out singleSwitchStates
		);
	end component singleSwitch_15;
	component singleSwitch_16 is
		port(
			clock : in std_logic;
			R13_command : in routeCommands;
			R52_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R56_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D07 : out singleSwitchStates
		);
	end component singleSwitch_16;
	component singleSwitch_17 is
		port(
			clock : in std_logic;
			R13_command : in routeCommands;
			R56_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D16 : out singleSwitchStates
		);
	end component singleSwitch_17;
	component singleSwitch_18 is
		port(
			clock : in std_logic;
			R4_command : in routeCommands;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			R72_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D19 : out singleSwitchStates
		);
	end component singleSwitch_18;
	component singleSwitch_19 is
		port(
			clock : in std_logic;
			R8_command : in routeCommands;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			R80_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D21 : out singleSwitchStates
		);
	end component singleSwitch_19;
	component singleSwitch_20 is
		port(
			clock : in std_logic;
			R16_command : in routeCommands;
			R60_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D24 : out singleSwitchStates
		);
	end component singleSwitch_20;
	component doubleSwitch is
		port(
			clock : in std_logic;
			indication : in dSwitch_type;
			command_in : in dSwitch_type;
			command_out : out dSwitch_type;
			correspondence : out dSwitch_type
		);
	end component doubleSwitch;
	component railwaySignal is
		port(
			clock : in std_logic;
			indication : in signal_type;
			command_in : in signal_type;
			command_out : out signal_type;
			correspondence : out signal_type
		);
	end component railwaySignal;
	component node_0 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R1_command : in routeCommands;
			R20_command : in routeCommands;
			R41_command : in routeCommands;
			R42_command : in routeCommands;
			R43_command : in routeCommands;
			R49_command : in routeCommands;
			state : out nodeStates
		);
	end component node_0;
	component node_1 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R37_command : in routeCommands;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			R58_command : in routeCommands;
			R69_command : in routeCommands;
			state : out nodeStates
		);
	end component node_1;
	component node_2 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			R36_command : in routeCommands;
			R38_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			state : out nodeStates
		);
	end component node_2;
	component node_3 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			state : out nodeStates
		);
	end component node_3;
	component node_4 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R40_command : in routeCommands;
			R59_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			R82_command : in routeCommands;
			state : out nodeStates
		);
	end component node_4;
	component node_5 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R26_command : in routeCommands;
			R28_command : in routeCommands;
			R39_command : in routeCommands;
			R80_command : in routeCommands;
			R81_command : in routeCommands;
			state : out nodeStates
		);
	end component node_5;
	component node_6 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R10_command : in routeCommands;
			R17_command : in routeCommands;
			R27_command : in routeCommands;
			R29_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			R78_command : in routeCommands;
			state : out nodeStates
		);
	end component node_6;
	component node_7 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R45_command : in routeCommands;
			R46_command : in routeCommands;
			R49_command : in routeCommands;
			state : out nodeStates
		);
	end component node_7;
	component node_8 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R2_command : in routeCommands;
			R20_command : in routeCommands;
			R22_command : in routeCommands;
			R42_command : in routeCommands;
			R66_command : in routeCommands;
			R67_command : in routeCommands;
			state : out nodeStates
		);
	end component node_8;
	component node_9 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R21_command : in routeCommands;
			R22_command : in routeCommands;
			R66_command : in routeCommands;
			R90_command : in routeCommands;
			state : out nodeStates
		);
	end component node_9;
	component node_10 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R43_command : in routeCommands;
			R45_command : in routeCommands;
			R47_command : in routeCommands;
			R50_command : in routeCommands;
			state : out nodeStates
		);
	end component node_10;
	component node_11 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R44_command : in routeCommands;
			R47_command : in routeCommands;
			R50_command : in routeCommands;
			R51_command : in routeCommands;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			R89_command : in routeCommands;
			R91_command : in routeCommands;
			state : out nodeStates
		);
	end component node_11;
	component node_12 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R2_command : in routeCommands;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			R67_command : in routeCommands;
			state : out nodeStates
		);
	end component node_12;
	component node_13 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R44_command : in routeCommands;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R51_command : in routeCommands;
			state : out nodeStates
		);
	end component node_13;
	component node_14 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R13_command : in routeCommands;
			R52_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R56_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			R65_command : in routeCommands;
			R86_command : in routeCommands;
			state : out nodeStates
		);
	end component node_14;
	component node_15 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R52_command : in routeCommands;
			R53_command : in routeCommands;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			state : out nodeStates
		);
	end component node_15;
	component node_16 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R13_command : in routeCommands;
			R54_command : in routeCommands;
			R56_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			state : out nodeStates
		);
	end component node_16;
	component node_17 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			R72_command : in routeCommands;
			state : out nodeStates
		);
	end component node_17;
	component node_18 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R7_command : in routeCommands;
			R77_command : in routeCommands;
			R79_command : in routeCommands;
			state : out nodeStates
		);
	end component node_18;
	component node_19 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			R80_command : in routeCommands;
			state : out nodeStates
		);
	end component node_19;
	component node_20 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R18_command : in routeCommands;
			R23_command : in routeCommands;
			R30_command : in routeCommands;
			R31_command : in routeCommands;
			R36_command : in routeCommands;
			R55_command : in routeCommands;
			R69_command : in routeCommands;
			state : out nodeStates
		);
	end component node_20;
	component node_21 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R30_command : in routeCommands;
			R36_command : in routeCommands;
			R37_command : in routeCommands;
			R38_command : in routeCommands;
			R55_command : in routeCommands;
			R69_command : in routeCommands;
			state : out nodeStates
		);
	end component node_21;
	component node_22 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R19_command : in routeCommands;
			R24_command : in routeCommands;
			R25_command : in routeCommands;
			R32_command : in routeCommands;
			R33_command : in routeCommands;
			R34_command : in routeCommands;
			R35_command : in routeCommands;
			state : out nodeStates
		);
	end component node_22;
	component node_23 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			R32_command : in routeCommands;
			R34_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			R59_command : in routeCommands;
			R82_command : in routeCommands;
			state : out nodeStates
		);
	end component node_23;
	component node_24 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R10_command : in routeCommands;
			R29_command : in routeCommands;
			state : out nodeStates
		);
	end component node_24;
	component node_25 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R48_command : in routeCommands;
			state : out nodeStates
		);
	end component node_25;
	component node_26 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R44_command : in routeCommands;
			R46_command : in routeCommands;
			R49_command : in routeCommands;
			state : out nodeStates
		);
	end component node_26;
	component node_27 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R2_command : in routeCommands;
			R67_command : in routeCommands;
			state : out nodeStates
		);
	end component node_27;
	component node_28 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			state : out nodeStates
		);
	end component node_28;
	component node_29 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R13_command : in routeCommands;
			R68_command : in routeCommands;
			state : out nodeStates
		);
	end component node_29;
	component node_30 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R69_command : in routeCommands;
			state : out nodeStates
		);
	end component node_30;
	component node_31 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			R72_command : in routeCommands;
			state : out nodeStates
		);
	end component node_31;
	component node_32 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			state : out nodeStates
		);
	end component node_32;
	component node_33 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R16_command : in routeCommands;
			R60_command : in routeCommands;
			R74_command : in routeCommands;
			R76_command : in routeCommands;
			R77_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			state : out nodeStates
		);
	end component node_33;
	component node_34 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			R78_command : in routeCommands;
			state : out nodeStates
		);
	end component node_34;
	component node_35 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R7_command : in routeCommands;
			R59_command : in routeCommands;
			R61_command : in routeCommands;
			R75_command : in routeCommands;
			R78_command : in routeCommands;
			R79_command : in routeCommands;
			state : out nodeStates
		);
	end component node_35;
	component node_36 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R80_command : in routeCommands;
			state : out nodeStates
		);
	end component node_36;
	component node_37 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R27_command : in routeCommands;
			R28_command : in routeCommands;
			R73_command : in routeCommands;
			R81_command : in routeCommands;
			state : out nodeStates
		);
	end component node_37;
	component node_38 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			state : out nodeStates
		);
	end component node_38;
	component node_39 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R16_command : in routeCommands;
			R83_command : in routeCommands;
			state : out nodeStates
		);
	end component node_39;
	component node_40 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R60_command : in routeCommands;
			R62_command : in routeCommands;
			R82_command : in routeCommands;
			state : out nodeStates
		);
	end component node_40;
	component node_41 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R24_command : in routeCommands;
			R33_command : in routeCommands;
			R65_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			state : out nodeStates
		);
	end component node_41;
	component node_42 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			state : out nodeStates
		);
	end component node_42;
	component node_43 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R65_command : in routeCommands;
			R86_command : in routeCommands;
			state : out nodeStates
		);
	end component node_43;
	component node_44 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			state : out nodeStates
		);
	end component node_44;
	component node_45 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R21_command : in routeCommands;
			R23_command : in routeCommands;
			R31_command : in routeCommands;
			R89_command : in routeCommands;
			R90_command : in routeCommands;
			R91_command : in routeCommands;
			state : out nodeStates
		);
	end component node_45;
	component node_46 is
		port(
			clock : in std_logic;
			ocupation : in std_logic;
			R89_command : in routeCommands;
			R91_command : in routeCommands;
			state : out nodeStates
		);
	end component node_46;
	component route_0 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne991_state : in nodeStates;
			ne991_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_0;
	component route_1 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne377_state : in nodeStates;
			ne377_command : out routeCommands;
			ne111_state : in nodeStates;
			ne111_command : out routeCommands;
			ne290_state : in nodeStates;
			ne290_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_1;
	component route_2 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne377_state : in nodeStates;
			ne377_command : out routeCommands;
			ne113_state : in nodeStates;
			ne113_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_2;
	component route_3 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne421_state : in nodeStates;
			ne421_command : out routeCommands;
			ne124_state : in nodeStates;
			ne124_command : out routeCommands;
			ne63_state : in nodeStates;
			ne63_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_3;
	component route_4 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne421_state : in nodeStates;
			ne421_command : out routeCommands;
			ne126_state : in nodeStates;
			ne126_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_4;
	component route_5 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne450_state : in nodeStates;
			ne450_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_5;
	component route_6 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne450_state : in nodeStates;
			ne450_command : out routeCommands;
			ne130_state : in nodeStates;
			ne130_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_6;
	component route_7 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne465_state : in nodeStates;
			ne465_command : out routeCommands;
			ne131_state : in nodeStates;
			ne131_command : out routeCommands;
			ne912_state : in nodeStates;
			ne912_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_7;
	component route_8 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne465_state : in nodeStates;
			ne465_command : out routeCommands;
			ne133_state : in nodeStates;
			ne133_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_8;
	component route_9 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne102_state : in nodeStates;
			ne102_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_9;
	component route_10 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne104_state : in nodeStates;
			ne104_command : out routeCommands;
			ne384_state : in nodeStates;
			ne384_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_10;
	component route_11 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne113_state : in nodeStates;
			ne113_command : out routeCommands;
			ne377_state : in nodeStates;
			ne377_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_11;
	component route_12 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne122_state : in nodeStates;
			ne122_command : out routeCommands;
			ne407_state : in nodeStates;
			ne407_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_12;
	component route_13 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne126_state : in nodeStates;
			ne126_command : out routeCommands;
			ne421_state : in nodeStates;
			ne421_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_13;
	component route_14 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne133_state : in nodeStates;
			ne133_command : out routeCommands;
			ne465_state : in nodeStates;
			ne465_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_14;
	component route_15 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne134_state : in nodeStates;
			ne134_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_15;
	component route_16 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_16;
	component route_17 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_17;
	component route_18 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_18;
	component route_19 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne290_state : in nodeStates;
			ne290_command : out routeCommands;
			ne991_state : in nodeStates;
			ne991_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_19;
	component route_20 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne292_state : in nodeStates;
			ne292_command : out routeCommands;
			ne996_state : in nodeStates;
			ne996_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_20;
	component route_21 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne292_state : in nodeStates;
			ne292_command : out routeCommands;
			ne290_state : in nodeStates;
			ne290_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_21;
	component route_22 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne996_state : in nodeStates;
			ne996_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_22;
	component route_23 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne992_state : in nodeStates;
			ne992_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_23;
	component route_24 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_24;
	component route_25 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne912_state : in nodeStates;
			ne912_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_25;
	component route_26 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne132_state : in nodeStates;
			ne132_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_26;
	component route_27 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne132_state : in nodeStates;
			ne132_command : out routeCommands;
			ne912_state : in nodeStates;
			ne912_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_27;
	component route_28 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			ne102_state : in nodeStates;
			ne102_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_28;
	component route_29 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_command : out routeCommands;
			Lc01_state : in levelCrossingStates;
			Lc01_command : out routeCommands;
			Lc02_state : in levelCrossingStates;
			Lc02_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_29;
	component route_30 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			ne996_state : in nodeStates;
			ne996_command : out routeCommands;
			Lc01_state : in levelCrossingStates;
			Lc01_command : out routeCommands;
			Lc02_state : in levelCrossingStates;
			Lc02_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_30;
	component route_31 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			Lc03_state : in levelCrossingStates;
			Lc03_command : out routeCommands;
			Lc04_state : in levelCrossingStates;
			Lc04_command : out routeCommands;
			Lc05_state : in levelCrossingStates;
			Lc05_command : out routeCommands;
			Lc06_state : in levelCrossingStates;
			Lc06_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_31;
	component route_32 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_command : out routeCommands;
			ne992_state : in nodeStates;
			ne992_command : out routeCommands;
			Lc03_state : in levelCrossingStates;
			Lc03_command : out routeCommands;
			Lc05_state : in levelCrossingStates;
			Lc05_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_32;
	component route_33 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			Lc04_state : in levelCrossingStates;
			Lc04_command : out routeCommands;
			Lc06_state : in levelCrossingStates;
			Lc06_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_33;
	component route_34 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_command : out routeCommands;
			Lc04_state : in levelCrossingStates;
			Lc04_command : out routeCommands;
			Lc06_state : in levelCrossingStates;
			Lc06_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_34;
	component route_35 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne63_state : in nodeStates;
			ne63_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_35;
	component route_36 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne99_state : in nodeStates;
			ne99_command : out routeCommands;
			ne61_state : in nodeStates;
			ne61_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_36;
	component route_37 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne99_state : in nodeStates;
			ne99_command : out routeCommands;
			ne63_state : in nodeStates;
			ne63_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_37;
	component route_38 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			ne912_state : in nodeStates;
			ne912_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_38;
	component route_39 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			ne910_state : in nodeStates;
			ne910_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_39;
	component route_40 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne991_state : in nodeStates;
			ne991_command : out routeCommands;
			ne288_state : in nodeStates;
			ne288_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_40;
	component route_41 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne991_state : in nodeStates;
			ne991_command : out routeCommands;
			ne290_state : in nodeStates;
			ne290_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_41;
	component route_42 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne295_state : in nodeStates;
			ne295_command : out routeCommands;
			ne288_state : in nodeStates;
			ne288_command : out routeCommands;
			ne991_state : in nodeStates;
			ne991_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_42;
	component route_43 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne110_state : in nodeStates;
			ne110_command : out routeCommands;
			ne384_state : in nodeStates;
			ne384_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_43;
	component route_44 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne288_state : in nodeStates;
			ne288_command : out routeCommands;
			ne295_state : in nodeStates;
			ne295_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_44;
	component route_45 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne288_state : in nodeStates;
			ne288_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_45;
	component route_46 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne295_state : in nodeStates;
			ne295_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_46;
	component route_47 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne384_state : in nodeStates;
			ne384_command : out routeCommands;
			ne104_state : in nodeStates;
			ne104_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_47;
	component route_48 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne384_state : in nodeStates;
			ne384_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_command : out routeCommands;
			ne288_state : in nodeStates;
			ne288_command : out routeCommands;
			ne991_state : in nodeStates;
			ne991_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_48;
	component route_49 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			ne295_state : in nodeStates;
			ne295_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_49;
	component route_50 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			ne384_state : in nodeStates;
			ne384_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_50;
	component route_51 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne404_state : in nodeStates;
			ne404_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_51;
	component route_52 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			ne404_state : in nodeStates;
			ne404_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_52;
	component route_53 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			ne407_state : in nodeStates;
			ne407_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_53;
	component route_54 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne404_state : in nodeStates;
			ne404_command : out routeCommands;
			ne61_state : in nodeStates;
			ne61_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_54;
	component route_55 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne123_state : in nodeStates;
			ne123_command : out routeCommands;
			ne407_state : in nodeStates;
			ne407_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_55;
	component route_56 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne61_state : in nodeStates;
			ne61_command : out routeCommands;
			ne404_state : in nodeStates;
			ne404_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_56;
	component route_57 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne61_state : in nodeStates;
			ne61_command : out routeCommands;
			ne123_state : in nodeStates;
			ne123_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_57;
	component route_58 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne130_state : in nodeStates;
			ne130_command : out routeCommands;
			ne910_state : in nodeStates;
			ne910_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_58;
	component route_59 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne135_state : in nodeStates;
			ne135_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_59;
	component route_60 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne910_state : in nodeStates;
			ne910_command : out routeCommands;
			ne130_state : in nodeStates;
			ne130_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_60;
	component route_61 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne910_state : in nodeStates;
			ne910_command : out routeCommands;
			ne135_state : in nodeStates;
			ne135_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_61;
	component route_62 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne993_state : in nodeStates;
			ne993_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_62;
	component route_63 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			ne993_state : in nodeStates;
			ne993_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_63;
	component route_64 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			ne994_state : in nodeStates;
			ne994_command : out routeCommands;
			ne992_state : in nodeStates;
			ne992_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_64;
	component route_65 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne290_state : in nodeStates;
			ne290_command : out routeCommands;
			ne292_state : in nodeStates;
			ne292_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_65;
	component route_66 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne290_state : in nodeStates;
			ne290_command : out routeCommands;
			ne111_state : in nodeStates;
			ne111_command : out routeCommands;
			ne377_state : in nodeStates;
			ne377_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_66;
	component route_67 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne407_state : in nodeStates;
			ne407_command : out routeCommands;
			ne122_state : in nodeStates;
			ne122_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_67;
	component route_68 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne407_state : in nodeStates;
			ne407_command : out routeCommands;
			ne123_state : in nodeStates;
			ne123_command : out routeCommands;
			ne61_state : in nodeStates;
			ne61_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_68;
	component route_69 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne65_state : in nodeStates;
			ne65_command : out routeCommands;
			ne63_state : in nodeStates;
			ne63_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_69;
	component route_70 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne63_state : in nodeStates;
			ne63_command : out routeCommands;
			ne65_state : in nodeStates;
			ne65_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_70;
	component route_71 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne63_state : in nodeStates;
			ne63_command : out routeCommands;
			ne124_state : in nodeStates;
			ne124_command : out routeCommands;
			ne421_state : in nodeStates;
			ne421_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_71;
	component route_72 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			ne132_state : in nodeStates;
			ne132_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_72;
	component route_73 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_73;
	component route_74 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_command : out routeCommands;
			ne130_state : in nodeStates;
			ne130_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_74;
	component route_75 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_75;
	component route_76 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			ne450_state : in nodeStates;
			ne450_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_76;
	component route_77 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne130_state : in nodeStates;
			ne130_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_77;
	component route_78 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne130_state : in nodeStates;
			ne130_command : out routeCommands;
			ne450_state : in nodeStates;
			ne450_command : out routeCommands;
			D12__state : in singleSwitchStates;
			D12__command : out routeCommands;
			routeState : out std_logic
		);
	end component route_78;
	component route_79 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne912_state : in nodeStates;
			ne912_command : out routeCommands;
			ne131_state : in nodeStates;
			ne131_command : out routeCommands;
			ne465_state : in nodeStates;
			ne465_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_79;
	component route_80 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne912_state : in nodeStates;
			ne912_command : out routeCommands;
			ne132_state : in nodeStates;
			ne132_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_80;
	component route_81 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			ne135_state : in nodeStates;
			ne135_command : out routeCommands;
			ne910_state : in nodeStates;
			ne910_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_81;
	component route_82 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_command : out routeCommands;
			ne134_state : in nodeStates;
			ne134_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_82;
	component route_83 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne65_state : in nodeStates;
			ne65_command : out routeCommands;
			ne992_state : in nodeStates;
			ne992_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_83;
	component route_84 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne992_state : in nodeStates;
			ne992_command : out routeCommands;
			ne65_state : in nodeStates;
			ne65_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_84;
	component route_85 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne992_state : in nodeStates;
			ne992_command : out routeCommands;
			ne994_state : in nodeStates;
			ne994_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_85;
	component route_86 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne995_state : in nodeStates;
			ne995_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_86;
	component route_87 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			ne995_state : in nodeStates;
			ne995_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_87;
	component route_88 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			ne997_state : in nodeStates;
			ne997_command : out routeCommands;
			ne996_state : in nodeStates;
			ne996_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_88;
	component route_89 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne996_state : in nodeStates;
			ne996_command : out routeCommands;
			ne292_state : in nodeStates;
			ne292_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_89;
	component route_90 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne996_state : in nodeStates;
			ne996_command : out routeCommands;
			ne997_state : in nodeStates;
			ne997_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_command : out routeCommands;
			routeState : out std_logic
		);
	end component route_90;

 signal state_Lc01 , state_Lc02 , state_Lc03 , state_Lc04 , state_Lc05 , state_Lc06 : levelCrossingStates;
 signal state_D01 , state_D08 , state_D05 , state_D18 , state_Sw01 , state_D10 , state_D09 , state_D20 , state_D23 , state_D03 , state_D14 , state_Sw04 , state_D04 , state_Sw03 , state_D15 , state_Sw02 , state_D07 , state_D16 , state_D19 , state_D21 , state_D24 : singleSwitchStates;
 signal state_ne991 , state_ne61 , state_ne63 , state_ne65 , state_ne910 , state_ne912 , state_ne114 , state_ne288 , state_ne290 , state_ne292 , state_ne295 , state_ne297 , state_ne377 , state_ne384 , state_ne400 , state_ne404 , state_ne407 , state_ne421 , state_ne450 , state_ne465 , state_ne98 , state_ne99 , state_ne100 , state_ne101 , state_ne102 , state_ne104 , state_ne110 , state_ne111 , state_ne113 , state_ne122 , state_ne123 , state_ne124 , state_ne126 , state_ne127 , state_ne129 , state_ne130 , state_ne131 , state_ne132 , state_ne133 , state_ne134 , state_ne135 , state_ne992 , state_ne993 , state_ne994 , state_ne995 , state_ne996 , state_ne997 : nodeStates;
 signal cmd_R1_ne991 , cmd_R2_ne377 , cmd_R2_ne111 , cmd_R2_ne290 , cmd_R3_ne377 , cmd_R3_ne113 , cmd_R4_ne421 , cmd_R4_ne124 , cmd_R4_ne63 , cmd_R5_ne421 , cmd_R5_ne126 , cmd_R6_ne450 , cmd_R6_ne127 , cmd_R7_ne450 , cmd_R7_ne130 , cmd_R8_ne465 , cmd_R8_ne131 , cmd_R8_ne912 , cmd_R9_ne465 , cmd_R9_ne133 , cmd_R10_ne102 , cmd_R10_ne114 , cmd_R11_ne104 , cmd_R11_ne384 , cmd_R11_ne297 , cmd_R12_ne113 , cmd_R12_ne377 , cmd_R13_ne122 , cmd_R13_ne407 , cmd_R13_ne400 , cmd_R14_ne126 , cmd_R14_ne421 , cmd_R15_ne133 , cmd_R15_ne465 , cmd_R16_ne134 , cmd_R16_ne127 , cmd_R17_ne114 , cmd_R18_ne98 , cmd_R19_ne100 , cmd_R20_ne290 , cmd_R20_ne991 , cmd_R21_ne292 , cmd_R21_ne996 , cmd_R22_ne292 , cmd_R22_ne290 , cmd_R23_ne996 , cmd_R23_ne98 , cmd_R24_ne992 , cmd_R24_ne100 , cmd_R25_ne101 , cmd_R25_ne100 , cmd_R26_ne912 , cmd_R26_ne101 , cmd_R27_ne132 , cmd_R27_ne114 , cmd_R28_ne132 , cmd_R28_ne912 , cmd_R29_ne114 , cmd_R29_ne102 , cmd_R30_ne98 , cmd_R30_ne99 , cmd_R31_ne98 , cmd_R31_ne996 , cmd_R32_ne100 , cmd_R32_ne101 , cmd_R33_ne100 , cmd_R33_ne992 , cmd_R34_ne100 , cmd_R34_ne101 , cmd_R35_ne100 , cmd_R36_ne63 , cmd_R36_ne99 , cmd_R36_ne98 , cmd_R37_ne99 , cmd_R37_ne61 , cmd_R38_ne99 , cmd_R38_ne63 , cmd_R39_ne101 , cmd_R39_ne912 , cmd_R40_ne101 , cmd_R40_ne910 , cmd_R41_ne991 , cmd_R41_ne288 , cmd_R42_ne991 , cmd_R42_ne290 , cmd_R43_ne295 , cmd_R43_ne288 , cmd_R43_ne991 , cmd_R44_ne110 , cmd_R44_ne384 , cmd_R44_ne297 , cmd_R45_ne288 , cmd_R45_ne295 , cmd_R46_ne288 , cmd_R46_ne110 , cmd_R47_ne295 , cmd_R47_ne297 , cmd_R48_ne384 , cmd_R48_ne104 , cmd_R49_ne384 , cmd_R49_ne110 , cmd_R49_ne288 , cmd_R49_ne991 , cmd_R50_ne297 , cmd_R50_ne295 , cmd_R51_ne297 , cmd_R51_ne384 , cmd_R52_ne404 , cmd_R52_ne400 , cmd_R53_ne400 , cmd_R53_ne404 , cmd_R54_ne400 , cmd_R54_ne407 , cmd_R55_ne404 , cmd_R55_ne61 , cmd_R55_ne99 , cmd_R55_ne98 , cmd_R56_ne123 , cmd_R56_ne407 , cmd_R56_ne400 , cmd_R57_ne61 , cmd_R57_ne404 , cmd_R58_ne61 , cmd_R58_ne123 , cmd_R59_ne130 , cmd_R59_ne910 , cmd_R59_ne101 , cmd_R60_ne135 , cmd_R60_ne127 , cmd_R61_ne910 , cmd_R61_ne130 , cmd_R62_ne910 , cmd_R62_ne135 , cmd_R63_ne993 , cmd_R63_ne400 , cmd_R64_ne400 , cmd_R64_ne993 , cmd_R65_ne400 , cmd_R65_ne994 , cmd_R65_ne992 , cmd_R66_ne290 , cmd_R66_ne292 , cmd_R67_ne290 , cmd_R67_ne111 , cmd_R67_ne377 , cmd_R68_ne407 , cmd_R68_ne122 , cmd_R69_ne407 , cmd_R69_ne123 , cmd_R69_ne61 , cmd_R69_ne99 , cmd_R69_ne98 , cmd_R70_ne65 , cmd_R70_ne63 , cmd_R71_ne63 , cmd_R71_ne65 , cmd_R72_ne63 , cmd_R72_ne124 , cmd_R72_ne421 , cmd_R73_ne114 , cmd_R73_ne132 , cmd_R74_ne114 , cmd_R74_ne129 , cmd_R74_ne127 , cmd_R75_ne114 , cmd_R75_ne129 , cmd_R75_ne130 , cmd_R76_ne127 , cmd_R76_ne129 , cmd_R76_ne114 , cmd_R77_ne127 , cmd_R77_ne450 , cmd_R78_ne130 , cmd_R78_ne129 , cmd_R78_ne114 , cmd_R79_ne130 , cmd_R79_ne450 , cmd_R80_ne912 , cmd_R80_ne131 , cmd_R80_ne465 , cmd_R81_ne912 , cmd_R81_ne132 , cmd_R82_ne127 , cmd_R82_ne135 , cmd_R82_ne910 , cmd_R82_ne101 , cmd_R83_ne127 , cmd_R83_ne134 , cmd_R84_ne65 , cmd_R84_ne992 , cmd_R85_ne992 , cmd_R85_ne65 , cmd_R86_ne992 , cmd_R86_ne994 , cmd_R86_ne400 , cmd_R87_ne995 , cmd_R87_ne297 , cmd_R88_ne297 , cmd_R88_ne995 , cmd_R89_ne297 , cmd_R89_ne997 , cmd_R89_ne996 , cmd_R90_ne996 , cmd_R90_ne292 , cmd_R91_ne996 , cmd_R91_ne997 , cmd_R91_ne297 : routeCommands;
 signal cmd_R30_Lc01 , cmd_R30_Lc02 , cmd_R31_Lc01 , cmd_R31_Lc02 , cmd_R32_Lc03 , cmd_R32_Lc04 , cmd_R32_Lc05 , cmd_R32_Lc06 , cmd_R33_Lc03 , cmd_R33_Lc05 , cmd_R34_Lc04 , cmd_R34_Lc06 , cmd_R35_Lc04 , cmd_R35_Lc06 : routeCommands;
 signal cmd_R2_D14 , cmd_R2_D15 , cmd_R3_D15 , cmd_R4_D18 , cmd_R4_D19 , cmd_R5_D19 , cmd_R6_D12_ , cmd_R7_D12_ , cmd_R8_D20 , cmd_R8_D21 , cmd_R9_D21 , cmd_R11_D04 , cmd_R12_D15 , cmd_R13_D07 , cmd_R13_D16 , cmd_R14_D19 , cmd_R15_D21 , cmd_R16_D24 , cmd_R20_D01 , cmd_R21_Sw04 , cmd_R22_D14 , cmd_R26_D09 , cmd_R27_D23 , cmd_R28_D20 , cmd_R36_D05 , cmd_R37_D05 , cmd_R38_D05 , cmd_R39_D09 , cmd_R40_D09 , cmd_R41_D01 , cmd_R42_D01 , cmd_R43_D01 , cmd_R43_D03 , cmd_R44_D04 , cmd_R45_D03 , cmd_R46_D03 , cmd_R47_D04 , cmd_R49_D01 , cmd_R49_D03 , cmd_R50_D04 , cmd_R51_D04 , cmd_R52_D07 , cmd_R53_D07 , cmd_R54_D07 , cmd_R55_D05 , cmd_R55_D08 , cmd_R56_D07 , cmd_R56_D16 , cmd_R57_D08 , cmd_R58_D08 , cmd_R59_D09 , cmd_R59_D10 , cmd_R60_D24 , cmd_R61_D10 , cmd_R62_D10 , cmd_R63_Sw02 , cmd_R64_Sw02 , cmd_R65_Sw02 , cmd_R65_Sw01 , cmd_R66_D14 , cmd_R67_D14 , cmd_R67_D15 , cmd_R68_D16 , cmd_R69_D05 , cmd_R69_D08 , cmd_R69_D16 , cmd_R70_D18 , cmd_R71_D18 , cmd_R72_D18 , cmd_R72_D19 , cmd_R73_D23 , cmd_R74_D23 , cmd_R74_D12_ , cmd_R75_D23 , cmd_R75_D12_ , cmd_R76_D23 , cmd_R76_D12_ , cmd_R77_D12_ , cmd_R78_D23 , cmd_R78_D12_ , cmd_R79_D12_ , cmd_R80_D20 , cmd_R80_D21 , cmd_R81_D20 , cmd_R82_D09 , cmd_R82_D10 , cmd_R82_D24 , cmd_R83_D24 , cmd_R84_Sw01 , cmd_R85_Sw01 , cmd_R86_Sw02 , cmd_R86_Sw01 , cmd_R87_Sw03 , cmd_R88_Sw03 , cmd_R89_Sw03 , cmd_R89_Sw04 , cmd_R90_Sw04 , cmd_R91_Sw03 , cmd_R91_Sw04 : routeCommands;
begin
	levelCrossing_Lc01 : levelCrossing_0 port map(clock => clock, R30_command => cmd_R30_Lc01, R31_command => cmd_R31_Lc01, ocupation_ne98 => ocupation(20), ocupation_ne996 => ocupation(45), ocupation_ne99 => ocupation(21), indication => levelCrossings_i(0), command  => levelCrossings_o(0), correspondence_Lc01 => state_Lc01);
	levelCrossing_Lc02 : levelCrossing_1 port map(clock => clock, R30_command => cmd_R30_Lc02, R31_command => cmd_R31_Lc02, ocupation_ne98 => ocupation(20), ocupation_ne996 => ocupation(45), ocupation_ne99 => ocupation(21), indication => levelCrossings_i(1), command  => levelCrossings_o(1), correspondence_Lc02 => state_Lc02);
	levelCrossing_Lc03 : levelCrossing_2 port map(clock => clock, R32_command => cmd_R32_Lc03, R33_command => cmd_R33_Lc03, ocupation_ne100 => ocupation(22), ocupation_ne992 => ocupation(41), ocupation_ne101 => ocupation(23), indication => levelCrossings_i(2), command  => levelCrossings_o(2), correspondence_Lc03 => state_Lc03);
	levelCrossing_Lc04 : levelCrossing_3 port map(clock => clock, R32_command => cmd_R32_Lc04, R34_command => cmd_R34_Lc04, R35_command => cmd_R35_Lc04, ocupation_ne100 => ocupation(22), ocupation_ne992 => ocupation(41), ocupation_ne101 => ocupation(23), indication => levelCrossings_i(3), command  => levelCrossings_o(3), correspondence_Lc04 => state_Lc04);
	levelCrossing_Lc05 : levelCrossing_4 port map(clock => clock, R32_command => cmd_R32_Lc05, R33_command => cmd_R33_Lc05, ocupation_ne100 => ocupation(22), ocupation_ne992 => ocupation(41), ocupation_ne101 => ocupation(23), indication => levelCrossings_i(4), command  => levelCrossings_o(4), correspondence_Lc05 => state_Lc05);
	levelCrossing_Lc06 : levelCrossing_5 port map(clock => clock, R32_command => cmd_R32_Lc06, R34_command => cmd_R34_Lc06, R35_command => cmd_R35_Lc06, ocupation_ne100 => ocupation(22), ocupation_ne992 => ocupation(41), ocupation_ne101 => ocupation(23), indication => levelCrossings_i(5), command  => levelCrossings_o(5), correspondence_Lc06 => state_Lc06);
	singleSwitch_D01 : singleSwitch_0 port map(clock => clock, R20_command => cmd_R20_D01, R41_command => cmd_R41_D01, R42_command => cmd_R42_D01, R43_command => cmd_R43_D01, R49_command => cmd_R49_D01, indication => singleSwitches_i(0), command => singleSwitches_o(0), correspondence_D01 => state_D01);
	singleSwitch_D08 : singleSwitch_1 port map(clock => clock, R55_command => cmd_R55_D08, R57_command => cmd_R57_D08, R58_command => cmd_R58_D08, R69_command => cmd_R69_D08, indication => singleSwitches_i(1), command => singleSwitches_o(1), correspondence_D08 => state_D08);
	singleSwitch_D05 : singleSwitch_2 port map(clock => clock, R36_command => cmd_R36_D05, R37_command => cmd_R37_D05, R38_command => cmd_R38_D05, R55_command => cmd_R55_D05, R69_command => cmd_R69_D05, indication => singleSwitches_i(2), command => singleSwitches_o(2), correspondence_D05 => state_D05);
	singleSwitch_D18 : singleSwitch_3 port map(clock => clock, R4_command => cmd_R4_D18, R70_command => cmd_R70_D18, R71_command => cmd_R71_D18, R72_command => cmd_R72_D18, indication => singleSwitches_i(3), command => singleSwitches_o(3), correspondence_D18 => state_D18);
	singleSwitch_Sw01 : singleSwitch_4 port map(clock => clock, R65_command => cmd_R65_Sw01, R84_command => cmd_R84_Sw01, R85_command => cmd_R85_Sw01, R86_command => cmd_R86_Sw01, indication => singleSwitches_i(4), command => singleSwitches_o(4), correspondence_Sw01 => state_Sw01);
	singleSwitch_D10 : singleSwitch_5 port map(clock => clock, R59_command => cmd_R59_D10, R61_command => cmd_R61_D10, R62_command => cmd_R62_D10, R82_command => cmd_R82_D10, indication => singleSwitches_i(5), command => singleSwitches_o(5), correspondence_D10 => state_D10);
	singleSwitch_D09 : singleSwitch_6 port map(clock => clock, R26_command => cmd_R26_D09, R39_command => cmd_R39_D09, R40_command => cmd_R40_D09, R59_command => cmd_R59_D09, R82_command => cmd_R82_D09, indication => singleSwitches_i(6), command => singleSwitches_o(6), correspondence_D09 => state_D09);
	singleSwitch_D20 : singleSwitch_7 port map(clock => clock, R8_command => cmd_R8_D20, R28_command => cmd_R28_D20, R80_command => cmd_R80_D20, R81_command => cmd_R81_D20, indication => singleSwitches_i(7), command => singleSwitches_o(7), correspondence_D20 => state_D20);
	singleSwitch_D23 : singleSwitch_8 port map(clock => clock, R27_command => cmd_R27_D23, R73_command => cmd_R73_D23, R74_command => cmd_R74_D23, R75_command => cmd_R75_D23, R76_command => cmd_R76_D23, R78_command => cmd_R78_D23, indication => singleSwitches_i(8), command => singleSwitches_o(8), correspondence_D23 => state_D23);
	singleSwitch_D03 : singleSwitch_9 port map(clock => clock, R43_command => cmd_R43_D03, R45_command => cmd_R45_D03, R46_command => cmd_R46_D03, R49_command => cmd_R49_D03, indication => singleSwitches_i(9), command => singleSwitches_o(9), correspondence_D03 => state_D03);
	singleSwitch_D14 : singleSwitch_10 port map(clock => clock, R2_command => cmd_R2_D14, R22_command => cmd_R22_D14, R66_command => cmd_R66_D14, R67_command => cmd_R67_D14, indication => singleSwitches_i(10), command => singleSwitches_o(10), correspondence_D14 => state_D14);
	singleSwitch_Sw04 : singleSwitch_11 port map(clock => clock, R21_command => cmd_R21_Sw04, R89_command => cmd_R89_Sw04, R90_command => cmd_R90_Sw04, R91_command => cmd_R91_Sw04, indication => singleSwitches_i(11), command => singleSwitches_o(11), correspondence_Sw04 => state_Sw04);
	singleSwitch_D04 : singleSwitch_12 port map(clock => clock, R11_command => cmd_R11_D04, R44_command => cmd_R44_D04, R47_command => cmd_R47_D04, R50_command => cmd_R50_D04, R51_command => cmd_R51_D04, indication => singleSwitches_i(12), command => singleSwitches_o(12), correspondence_D04 => state_D04);
	singleSwitch_Sw03 : singleSwitch_13 port map(clock => clock, R87_command => cmd_R87_Sw03, R88_command => cmd_R88_Sw03, R89_command => cmd_R89_Sw03, R91_command => cmd_R91_Sw03, indication => singleSwitches_i(13), command => singleSwitches_o(13), correspondence_Sw03 => state_Sw03);
	singleSwitch_D15 : singleSwitch_14 port map(clock => clock, R2_command => cmd_R2_D15, R3_command => cmd_R3_D15, R12_command => cmd_R12_D15, R67_command => cmd_R67_D15, indication => singleSwitches_i(14), command => singleSwitches_o(14), correspondence_D15 => state_D15);
	singleSwitch_Sw02 : singleSwitch_15 port map(clock => clock, R63_command => cmd_R63_Sw02, R64_command => cmd_R64_Sw02, R65_command => cmd_R65_Sw02, R86_command => cmd_R86_Sw02, indication => singleSwitches_i(15), command => singleSwitches_o(15), correspondence_Sw02 => state_Sw02);
	singleSwitch_D07 : singleSwitch_16 port map(clock => clock, R13_command => cmd_R13_D07, R52_command => cmd_R52_D07, R53_command => cmd_R53_D07, R54_command => cmd_R54_D07, R56_command => cmd_R56_D07, indication => singleSwitches_i(16), command => singleSwitches_o(16), correspondence_D07 => state_D07);
	singleSwitch_D16 : singleSwitch_17 port map(clock => clock, R13_command => cmd_R13_D16, R56_command => cmd_R56_D16, R68_command => cmd_R68_D16, R69_command => cmd_R69_D16, indication => singleSwitches_i(17), command => singleSwitches_o(17), correspondence_D16 => state_D16);
	singleSwitch_D19 : singleSwitch_18 port map(clock => clock, R4_command => cmd_R4_D19, R5_command => cmd_R5_D19, R14_command => cmd_R14_D19, R72_command => cmd_R72_D19, indication => singleSwitches_i(18), command => singleSwitches_o(18), correspondence_D19 => state_D19);
	singleSwitch_D21 : singleSwitch_19 port map(clock => clock, R8_command => cmd_R8_D21, R9_command => cmd_R9_D21, R15_command => cmd_R15_D21, R80_command => cmd_R80_D21, indication => singleSwitches_i(19), command => singleSwitches_o(19), correspondence_D21 => state_D21);
	singleSwitch_D24 : singleSwitch_20 port map(clock => clock, R16_command => cmd_R16_D24, R60_command => cmd_R60_D24, R82_command => cmd_R82_D24, R83_command => cmd_R83_D24, indication => singleSwitches_i(20), command => singleSwitches_o(20), correspondence_D24 => state_D24);
	node_ne991 : node_0 port map(clock => clock, ocupation => ocupation(0), R1_command => cmd_R1_ne991, R20_command => cmd_R20_ne991, R41_command => cmd_R41_ne991, R42_command => cmd_R42_ne991, R43_command => cmd_R43_ne991, R49_command => cmd_R49_ne991, state => state_ne991);
	node_ne61 : node_1 port map(clock => clock, ocupation => ocupation(1), R37_command => cmd_R37_ne61, R55_command => cmd_R55_ne61, R57_command => cmd_R57_ne61, R58_command => cmd_R58_ne61, R69_command => cmd_R69_ne61, state => state_ne61);
	node_ne63 : node_2 port map(clock => clock, ocupation => ocupation(2), R4_command => cmd_R4_ne63, R36_command => cmd_R36_ne63, R38_command => cmd_R38_ne63, R70_command => cmd_R70_ne63, R71_command => cmd_R71_ne63, R72_command => cmd_R72_ne63, state => state_ne63);
	node_ne65 : node_3 port map(clock => clock, ocupation => ocupation(3), R70_command => cmd_R70_ne65, R71_command => cmd_R71_ne65, R84_command => cmd_R84_ne65, R85_command => cmd_R85_ne65, state => state_ne65);
	node_ne910 : node_4 port map(clock => clock, ocupation => ocupation(4), R40_command => cmd_R40_ne910, R59_command => cmd_R59_ne910, R61_command => cmd_R61_ne910, R62_command => cmd_R62_ne910, R82_command => cmd_R82_ne910, state => state_ne910);
	node_ne912 : node_5 port map(clock => clock, ocupation => ocupation(5), R8_command => cmd_R8_ne912, R26_command => cmd_R26_ne912, R28_command => cmd_R28_ne912, R39_command => cmd_R39_ne912, R80_command => cmd_R80_ne912, R81_command => cmd_R81_ne912, state => state_ne912);
	node_ne114 : node_6 port map(clock => clock, ocupation => ocupation(6), R10_command => cmd_R10_ne114, R17_command => cmd_R17_ne114, R27_command => cmd_R27_ne114, R29_command => cmd_R29_ne114, R73_command => cmd_R73_ne114, R74_command => cmd_R74_ne114, R75_command => cmd_R75_ne114, R76_command => cmd_R76_ne114, R78_command => cmd_R78_ne114, state => state_ne114);
	node_ne288 : node_7 port map(clock => clock, ocupation => ocupation(7), R41_command => cmd_R41_ne288, R43_command => cmd_R43_ne288, R45_command => cmd_R45_ne288, R46_command => cmd_R46_ne288, R49_command => cmd_R49_ne288, state => state_ne288);
	node_ne290 : node_8 port map(clock => clock, ocupation => ocupation(8), R2_command => cmd_R2_ne290, R20_command => cmd_R20_ne290, R22_command => cmd_R22_ne290, R42_command => cmd_R42_ne290, R66_command => cmd_R66_ne290, R67_command => cmd_R67_ne290, state => state_ne290);
	node_ne292 : node_9 port map(clock => clock, ocupation => ocupation(9), R21_command => cmd_R21_ne292, R22_command => cmd_R22_ne292, R66_command => cmd_R66_ne292, R90_command => cmd_R90_ne292, state => state_ne292);
	node_ne295 : node_10 port map(clock => clock, ocupation => ocupation(10), R43_command => cmd_R43_ne295, R45_command => cmd_R45_ne295, R47_command => cmd_R47_ne295, R50_command => cmd_R50_ne295, state => state_ne295);
	node_ne297 : node_11 port map(clock => clock, ocupation => ocupation(11), R11_command => cmd_R11_ne297, R44_command => cmd_R44_ne297, R47_command => cmd_R47_ne297, R50_command => cmd_R50_ne297, R51_command => cmd_R51_ne297, R87_command => cmd_R87_ne297, R88_command => cmd_R88_ne297, R89_command => cmd_R89_ne297, R91_command => cmd_R91_ne297, state => state_ne297);
	node_ne377 : node_12 port map(clock => clock, ocupation => ocupation(12), R2_command => cmd_R2_ne377, R3_command => cmd_R3_ne377, R12_command => cmd_R12_ne377, R67_command => cmd_R67_ne377, state => state_ne377);
	node_ne384 : node_13 port map(clock => clock, ocupation => ocupation(13), R11_command => cmd_R11_ne384, R44_command => cmd_R44_ne384, R48_command => cmd_R48_ne384, R49_command => cmd_R49_ne384, R51_command => cmd_R51_ne384, state => state_ne384);
	node_ne400 : node_14 port map(clock => clock, ocupation => ocupation(14), R13_command => cmd_R13_ne400, R52_command => cmd_R52_ne400, R53_command => cmd_R53_ne400, R54_command => cmd_R54_ne400, R56_command => cmd_R56_ne400, R63_command => cmd_R63_ne400, R64_command => cmd_R64_ne400, R65_command => cmd_R65_ne400, R86_command => cmd_R86_ne400, state => state_ne400);
	node_ne404 : node_15 port map(clock => clock, ocupation => ocupation(15), R52_command => cmd_R52_ne404, R53_command => cmd_R53_ne404, R55_command => cmd_R55_ne404, R57_command => cmd_R57_ne404, state => state_ne404);
	node_ne407 : node_16 port map(clock => clock, ocupation => ocupation(16), R13_command => cmd_R13_ne407, R54_command => cmd_R54_ne407, R56_command => cmd_R56_ne407, R68_command => cmd_R68_ne407, R69_command => cmd_R69_ne407, state => state_ne407);
	node_ne421 : node_17 port map(clock => clock, ocupation => ocupation(17), R4_command => cmd_R4_ne421, R5_command => cmd_R5_ne421, R14_command => cmd_R14_ne421, R72_command => cmd_R72_ne421, state => state_ne421);
	node_ne450 : node_18 port map(clock => clock, ocupation => ocupation(18), R6_command => cmd_R6_ne450, R7_command => cmd_R7_ne450, R77_command => cmd_R77_ne450, R79_command => cmd_R79_ne450, state => state_ne450);
	node_ne465 : node_19 port map(clock => clock, ocupation => ocupation(19), R8_command => cmd_R8_ne465, R9_command => cmd_R9_ne465, R15_command => cmd_R15_ne465, R80_command => cmd_R80_ne465, state => state_ne465);
	node_ne98 : node_20 port map(clock => clock, ocupation => ocupation(20), R18_command => cmd_R18_ne98, R23_command => cmd_R23_ne98, R30_command => cmd_R30_ne98, R31_command => cmd_R31_ne98, R36_command => cmd_R36_ne98, R55_command => cmd_R55_ne98, R69_command => cmd_R69_ne98, state => state_ne98);
	node_ne99 : node_21 port map(clock => clock, ocupation => ocupation(21), R30_command => cmd_R30_ne99, R36_command => cmd_R36_ne99, R37_command => cmd_R37_ne99, R38_command => cmd_R38_ne99, R55_command => cmd_R55_ne99, R69_command => cmd_R69_ne99, state => state_ne99);
	node_ne100 : node_22 port map(clock => clock, ocupation => ocupation(22), R19_command => cmd_R19_ne100, R24_command => cmd_R24_ne100, R25_command => cmd_R25_ne100, R32_command => cmd_R32_ne100, R33_command => cmd_R33_ne100, R34_command => cmd_R34_ne100, R35_command => cmd_R35_ne100, state => state_ne100);
	node_ne101 : node_23 port map(clock => clock, ocupation => ocupation(23), R25_command => cmd_R25_ne101, R26_command => cmd_R26_ne101, R32_command => cmd_R32_ne101, R34_command => cmd_R34_ne101, R39_command => cmd_R39_ne101, R40_command => cmd_R40_ne101, R59_command => cmd_R59_ne101, R82_command => cmd_R82_ne101, state => state_ne101);
	node_ne102 : node_24 port map(clock => clock, ocupation => ocupation(24), R10_command => cmd_R10_ne102, R29_command => cmd_R29_ne102, state => state_ne102);
	node_ne104 : node_25 port map(clock => clock, ocupation => ocupation(25), R11_command => cmd_R11_ne104, R48_command => cmd_R48_ne104, state => state_ne104);
	node_ne110 : node_26 port map(clock => clock, ocupation => ocupation(26), R44_command => cmd_R44_ne110, R46_command => cmd_R46_ne110, R49_command => cmd_R49_ne110, state => state_ne110);
	node_ne111 : node_27 port map(clock => clock, ocupation => ocupation(27), R2_command => cmd_R2_ne111, R67_command => cmd_R67_ne111, state => state_ne111);
	node_ne113 : node_28 port map(clock => clock, ocupation => ocupation(28), R3_command => cmd_R3_ne113, R12_command => cmd_R12_ne113, state => state_ne113);
	node_ne122 : node_29 port map(clock => clock, ocupation => ocupation(29), R13_command => cmd_R13_ne122, R68_command => cmd_R68_ne122, state => state_ne122);
	node_ne123 : node_30 port map(clock => clock, ocupation => ocupation(30), R56_command => cmd_R56_ne123, R58_command => cmd_R58_ne123, R69_command => cmd_R69_ne123, state => state_ne123);
	node_ne124 : node_31 port map(clock => clock, ocupation => ocupation(31), R4_command => cmd_R4_ne124, R72_command => cmd_R72_ne124, state => state_ne124);
	node_ne126 : node_32 port map(clock => clock, ocupation => ocupation(32), R5_command => cmd_R5_ne126, R14_command => cmd_R14_ne126, state => state_ne126);
	node_ne127 : node_33 port map(clock => clock, ocupation => ocupation(33), R6_command => cmd_R6_ne127, R16_command => cmd_R16_ne127, R60_command => cmd_R60_ne127, R74_command => cmd_R74_ne127, R76_command => cmd_R76_ne127, R77_command => cmd_R77_ne127, R82_command => cmd_R82_ne127, R83_command => cmd_R83_ne127, state => state_ne127);
	node_ne129 : node_34 port map(clock => clock, ocupation => ocupation(34), R74_command => cmd_R74_ne129, R75_command => cmd_R75_ne129, R76_command => cmd_R76_ne129, R78_command => cmd_R78_ne129, state => state_ne129);
	node_ne130 : node_35 port map(clock => clock, ocupation => ocupation(35), R7_command => cmd_R7_ne130, R59_command => cmd_R59_ne130, R61_command => cmd_R61_ne130, R75_command => cmd_R75_ne130, R78_command => cmd_R78_ne130, R79_command => cmd_R79_ne130, state => state_ne130);
	node_ne131 : node_36 port map(clock => clock, ocupation => ocupation(36), R8_command => cmd_R8_ne131, R80_command => cmd_R80_ne131, state => state_ne131);
	node_ne132 : node_37 port map(clock => clock, ocupation => ocupation(37), R27_command => cmd_R27_ne132, R28_command => cmd_R28_ne132, R73_command => cmd_R73_ne132, R81_command => cmd_R81_ne132, state => state_ne132);
	node_ne133 : node_38 port map(clock => clock, ocupation => ocupation(38), R9_command => cmd_R9_ne133, R15_command => cmd_R15_ne133, state => state_ne133);
	node_ne134 : node_39 port map(clock => clock, ocupation => ocupation(39), R16_command => cmd_R16_ne134, R83_command => cmd_R83_ne134, state => state_ne134);
	node_ne135 : node_40 port map(clock => clock, ocupation => ocupation(40), R60_command => cmd_R60_ne135, R62_command => cmd_R62_ne135, R82_command => cmd_R82_ne135, state => state_ne135);
	node_ne992 : node_41 port map(clock => clock, ocupation => ocupation(41), R24_command => cmd_R24_ne992, R33_command => cmd_R33_ne992, R65_command => cmd_R65_ne992, R84_command => cmd_R84_ne992, R85_command => cmd_R85_ne992, R86_command => cmd_R86_ne992, state => state_ne992);
	node_ne993 : node_42 port map(clock => clock, ocupation => ocupation(42), R63_command => cmd_R63_ne993, R64_command => cmd_R64_ne993, state => state_ne993);
	node_ne994 : node_43 port map(clock => clock, ocupation => ocupation(43), R65_command => cmd_R65_ne994, R86_command => cmd_R86_ne994, state => state_ne994);
	node_ne995 : node_44 port map(clock => clock, ocupation => ocupation(44), R87_command => cmd_R87_ne995, R88_command => cmd_R88_ne995, state => state_ne995);
	node_ne996 : node_45 port map(clock => clock, ocupation => ocupation(45), R21_command => cmd_R21_ne996, R23_command => cmd_R23_ne996, R31_command => cmd_R31_ne996, R89_command => cmd_R89_ne996, R90_command => cmd_R90_ne996, R91_command => cmd_R91_ne996, state => state_ne996);
	node_ne997 : node_46 port map(clock => clock, ocupation => ocupation(46), R89_command => cmd_R89_ne997, R91_command => cmd_R91_ne997, state => state_ne997);
	route_R1 : route_0 port map(clock => clock, routeRequest => routes_i(0), ne991_command => cmd_R1_ne991, ne991_state => state_ne991, routeState => routes_o(0));
	route_R2 : route_1 port map(clock => clock, routeRequest => routes_i(1), ne290_command => cmd_R2_ne290, ne290_state => state_ne290, ne377_command => cmd_R2_ne377, ne377_state => state_ne377, ne111_command => cmd_R2_ne111, ne111_state => state_ne111, D14_command => cmd_R2_D14, D14_state => state_D14, D15_command => cmd_R2_D15, D15_state => state_D15, routeState => routes_o(1));
	route_R3 : route_2 port map(clock => clock, routeRequest => routes_i(2), ne377_command => cmd_R3_ne377, ne377_state => state_ne377, ne113_command => cmd_R3_ne113, ne113_state => state_ne113, D15_command => cmd_R3_D15, D15_state => state_D15, routeState => routes_o(2));
	route_R4 : route_3 port map(clock => clock, routeRequest => routes_i(3), ne63_command => cmd_R4_ne63, ne63_state => state_ne63, ne421_command => cmd_R4_ne421, ne421_state => state_ne421, ne124_command => cmd_R4_ne124, ne124_state => state_ne124, D18_command => cmd_R4_D18, D18_state => state_D18, D19_command => cmd_R4_D19, D19_state => state_D19, routeState => routes_o(3));
	route_R5 : route_4 port map(clock => clock, routeRequest => routes_i(4), ne421_command => cmd_R5_ne421, ne421_state => state_ne421, ne126_command => cmd_R5_ne126, ne126_state => state_ne126, D19_command => cmd_R5_D19, D19_state => state_D19, routeState => routes_o(4));
	route_R6 : route_5 port map(clock => clock, routeRequest => routes_i(5), ne450_command => cmd_R6_ne450, ne450_state => state_ne450, ne127_command => cmd_R6_ne127, ne127_state => state_ne127, D12__command => cmd_R6_D12_, D12__state => state_D12_, routeState => routes_o(5));
	route_R7 : route_6 port map(clock => clock, routeRequest => routes_i(6), ne450_command => cmd_R7_ne450, ne450_state => state_ne450, ne130_command => cmd_R7_ne130, ne130_state => state_ne130, D12__command => cmd_R7_D12_, D12__state => state_D12_, routeState => routes_o(6));
	route_R8 : route_7 port map(clock => clock, routeRequest => routes_i(7), ne912_command => cmd_R8_ne912, ne912_state => state_ne912, ne465_command => cmd_R8_ne465, ne465_state => state_ne465, ne131_command => cmd_R8_ne131, ne131_state => state_ne131, D20_command => cmd_R8_D20, D20_state => state_D20, D21_command => cmd_R8_D21, D21_state => state_D21, routeState => routes_o(7));
	route_R9 : route_8 port map(clock => clock, routeRequest => routes_i(8), ne465_command => cmd_R9_ne465, ne465_state => state_ne465, ne133_command => cmd_R9_ne133, ne133_state => state_ne133, D21_command => cmd_R9_D21, D21_state => state_D21, routeState => routes_o(8));
	route_R10 : route_9 port map(clock => clock, routeRequest => routes_i(9), ne114_command => cmd_R10_ne114, ne114_state => state_ne114, ne102_command => cmd_R10_ne102, ne102_state => state_ne102, routeState => routes_o(9));
	route_R11 : route_10 port map(clock => clock, routeRequest => routes_i(10), ne297_command => cmd_R11_ne297, ne297_state => state_ne297, ne384_command => cmd_R11_ne384, ne384_state => state_ne384, ne104_command => cmd_R11_ne104, ne104_state => state_ne104, D04_command => cmd_R11_D04, D04_state => state_D04, routeState => routes_o(10));
	route_R12 : route_11 port map(clock => clock, routeRequest => routes_i(11), ne377_command => cmd_R12_ne377, ne377_state => state_ne377, ne113_command => cmd_R12_ne113, ne113_state => state_ne113, D15_command => cmd_R12_D15, D15_state => state_D15, routeState => routes_o(11));
	route_R13 : route_12 port map(clock => clock, routeRequest => routes_i(12), ne400_command => cmd_R13_ne400, ne400_state => state_ne400, ne407_command => cmd_R13_ne407, ne407_state => state_ne407, ne122_command => cmd_R13_ne122, ne122_state => state_ne122, D07_command => cmd_R13_D07, D07_state => state_D07, D16_command => cmd_R13_D16, D16_state => state_D16, routeState => routes_o(12));
	route_R14 : route_13 port map(clock => clock, routeRequest => routes_i(13), ne421_command => cmd_R14_ne421, ne421_state => state_ne421, ne126_command => cmd_R14_ne126, ne126_state => state_ne126, D19_command => cmd_R14_D19, D19_state => state_D19, routeState => routes_o(13));
	route_R15 : route_14 port map(clock => clock, routeRequest => routes_i(14), ne465_command => cmd_R15_ne465, ne465_state => state_ne465, ne133_command => cmd_R15_ne133, ne133_state => state_ne133, D21_command => cmd_R15_D21, D21_state => state_D21, routeState => routes_o(14));
	route_R16 : route_15 port map(clock => clock, routeRequest => routes_i(15), ne127_command => cmd_R16_ne127, ne127_state => state_ne127, ne134_command => cmd_R16_ne134, ne134_state => state_ne134, D24_command => cmd_R16_D24, D24_state => state_D24, routeState => routes_o(15));
	route_R17 : route_16 port map(clock => clock, routeRequest => routes_i(16), ne114_command => cmd_R17_ne114, ne114_state => state_ne114, routeState => routes_o(16));
	route_R18 : route_17 port map(clock => clock, routeRequest => routes_i(17), ne98_command => cmd_R18_ne98, ne98_state => state_ne98, routeState => routes_o(17));
	route_R19 : route_18 port map(clock => clock, routeRequest => routes_i(18), ne100_command => cmd_R19_ne100, ne100_state => state_ne100, routeState => routes_o(18));
	route_R20 : route_19 port map(clock => clock, routeRequest => routes_i(19), ne991_command => cmd_R20_ne991, ne991_state => state_ne991, ne290_command => cmd_R20_ne290, ne290_state => state_ne290, D01_command => cmd_R20_D01, D01_state => state_D01, routeState => routes_o(19));
	route_R21 : route_20 port map(clock => clock, routeRequest => routes_i(20), ne292_command => cmd_R21_ne292, ne292_state => state_ne292, ne996_command => cmd_R21_ne996, ne996_state => state_ne996, Sw04_command => cmd_R21_Sw04, Sw04_state => state_Sw04, routeState => routes_o(20));
	route_R22 : route_21 port map(clock => clock, routeRequest => routes_i(21), ne290_command => cmd_R22_ne290, ne290_state => state_ne290, ne292_command => cmd_R22_ne292, ne292_state => state_ne292, D14_command => cmd_R22_D14, D14_state => state_D14, routeState => routes_o(21));
	route_R23 : route_22 port map(clock => clock, routeRequest => routes_i(22), ne98_command => cmd_R23_ne98, ne98_state => state_ne98, ne996_command => cmd_R23_ne996, ne996_state => state_ne996, routeState => routes_o(22));
	route_R24 : route_23 port map(clock => clock, routeRequest => routes_i(23), ne100_command => cmd_R24_ne100, ne100_state => state_ne100, ne992_command => cmd_R24_ne992, ne992_state => state_ne992, routeState => routes_o(23));
	route_R25 : route_24 port map(clock => clock, routeRequest => routes_i(24), ne100_command => cmd_R25_ne100, ne100_state => state_ne100, ne101_command => cmd_R25_ne101, ne101_state => state_ne101, routeState => routes_o(24));
	route_R26 : route_25 port map(clock => clock, routeRequest => routes_i(25), ne912_command => cmd_R26_ne912, ne912_state => state_ne912, ne101_command => cmd_R26_ne101, ne101_state => state_ne101, D09_command => cmd_R26_D09, D09_state => state_D09, routeState => routes_o(25));
	route_R27 : route_26 port map(clock => clock, routeRequest => routes_i(26), ne114_command => cmd_R27_ne114, ne114_state => state_ne114, ne132_command => cmd_R27_ne132, ne132_state => state_ne132, D23_command => cmd_R27_D23, D23_state => state_D23, routeState => routes_o(26));
	route_R28 : route_27 port map(clock => clock, routeRequest => routes_i(27), ne912_command => cmd_R28_ne912, ne912_state => state_ne912, ne132_command => cmd_R28_ne132, ne132_state => state_ne132, D20_command => cmd_R28_D20, D20_state => state_D20, routeState => routes_o(27));
	route_R29 : route_28 port map(clock => clock, routeRequest => routes_i(28), ne114_command => cmd_R29_ne114, ne114_state => state_ne114, ne102_command => cmd_R29_ne102, ne102_state => state_ne102, routeState => routes_o(28));
	route_R30 : route_29 port map(clock => clock, routeRequest => routes_i(29), ne98_command => cmd_R30_ne98, ne98_state => state_ne98, ne99_command => cmd_R30_ne99, ne99_state => state_ne99, Lc01_command => cmd_R30_Lc01, Lc01_state => state_Lc01, Lc02_command => cmd_R30_Lc02, Lc02_state => state_Lc02, routeState => routes_o(29));
	route_R31 : route_30 port map(clock => clock, routeRequest => routes_i(30), ne98_command => cmd_R31_ne98, ne98_state => state_ne98, ne996_command => cmd_R31_ne996, ne996_state => state_ne996, Lc01_command => cmd_R31_Lc01, Lc01_state => state_Lc01, Lc02_command => cmd_R31_Lc02, Lc02_state => state_Lc02, routeState => routes_o(30));
	route_R32 : route_31 port map(clock => clock, routeRequest => routes_i(31), ne100_command => cmd_R32_ne100, ne100_state => state_ne100, ne101_command => cmd_R32_ne101, ne101_state => state_ne101, Lc03_command => cmd_R32_Lc03, Lc03_state => state_Lc03, Lc04_command => cmd_R32_Lc04, Lc04_state => state_Lc04, Lc05_command => cmd_R32_Lc05, Lc05_state => state_Lc05, Lc06_command => cmd_R32_Lc06, Lc06_state => state_Lc06, routeState => routes_o(31));
	route_R33 : route_32 port map(clock => clock, routeRequest => routes_i(32), ne100_command => cmd_R33_ne100, ne100_state => state_ne100, ne992_command => cmd_R33_ne992, ne992_state => state_ne992, Lc03_command => cmd_R33_Lc03, Lc03_state => state_Lc03, Lc05_command => cmd_R33_Lc05, Lc05_state => state_Lc05, routeState => routes_o(32));
	route_R34 : route_33 port map(clock => clock, routeRequest => routes_i(33), ne100_command => cmd_R34_ne100, ne100_state => state_ne100, ne101_command => cmd_R34_ne101, ne101_state => state_ne101, Lc04_command => cmd_R34_Lc04, Lc04_state => state_Lc04, Lc06_command => cmd_R34_Lc06, Lc06_state => state_Lc06, routeState => routes_o(33));
	route_R35 : route_34 port map(clock => clock, routeRequest => routes_i(34), ne100_command => cmd_R35_ne100, ne100_state => state_ne100, Lc04_command => cmd_R35_Lc04, Lc04_state => state_Lc04, Lc06_command => cmd_R35_Lc06, Lc06_state => state_Lc06, routeState => routes_o(34));
	route_R36 : route_35 port map(clock => clock, routeRequest => routes_i(35), ne63_command => cmd_R36_ne63, ne63_state => state_ne63, ne98_command => cmd_R36_ne98, ne98_state => state_ne98, ne99_command => cmd_R36_ne99, ne99_state => state_ne99, D05_command => cmd_R36_D05, D05_state => state_D05, routeState => routes_o(35));
	route_R37 : route_36 port map(clock => clock, routeRequest => routes_i(36), ne61_command => cmd_R37_ne61, ne61_state => state_ne61, ne99_command => cmd_R37_ne99, ne99_state => state_ne99, D05_command => cmd_R37_D05, D05_state => state_D05, routeState => routes_o(36));
	route_R38 : route_37 port map(clock => clock, routeRequest => routes_i(37), ne63_command => cmd_R38_ne63, ne63_state => state_ne63, ne99_command => cmd_R38_ne99, ne99_state => state_ne99, D05_command => cmd_R38_D05, D05_state => state_D05, routeState => routes_o(37));
	route_R39 : route_38 port map(clock => clock, routeRequest => routes_i(38), ne912_command => cmd_R39_ne912, ne912_state => state_ne912, ne101_command => cmd_R39_ne101, ne101_state => state_ne101, D09_command => cmd_R39_D09, D09_state => state_D09, routeState => routes_o(38));
	route_R40 : route_39 port map(clock => clock, routeRequest => routes_i(39), ne910_command => cmd_R40_ne910, ne910_state => state_ne910, ne101_command => cmd_R40_ne101, ne101_state => state_ne101, D09_command => cmd_R40_D09, D09_state => state_D09, routeState => routes_o(39));
	route_R41 : route_40 port map(clock => clock, routeRequest => routes_i(40), ne991_command => cmd_R41_ne991, ne991_state => state_ne991, ne288_command => cmd_R41_ne288, ne288_state => state_ne288, D01_command => cmd_R41_D01, D01_state => state_D01, routeState => routes_o(40));
	route_R42 : route_41 port map(clock => clock, routeRequest => routes_i(41), ne991_command => cmd_R42_ne991, ne991_state => state_ne991, ne290_command => cmd_R42_ne290, ne290_state => state_ne290, D01_command => cmd_R42_D01, D01_state => state_D01, routeState => routes_o(41));
	route_R43 : route_42 port map(clock => clock, routeRequest => routes_i(42), ne991_command => cmd_R43_ne991, ne991_state => state_ne991, ne288_command => cmd_R43_ne288, ne288_state => state_ne288, ne295_command => cmd_R43_ne295, ne295_state => state_ne295, D01_command => cmd_R43_D01, D01_state => state_D01, D03_command => cmd_R43_D03, D03_state => state_D03, routeState => routes_o(42));
	route_R44 : route_43 port map(clock => clock, routeRequest => routes_i(43), ne297_command => cmd_R44_ne297, ne297_state => state_ne297, ne384_command => cmd_R44_ne384, ne384_state => state_ne384, ne110_command => cmd_R44_ne110, ne110_state => state_ne110, D04_command => cmd_R44_D04, D04_state => state_D04, routeState => routes_o(43));
	route_R45 : route_44 port map(clock => clock, routeRequest => routes_i(44), ne288_command => cmd_R45_ne288, ne288_state => state_ne288, ne295_command => cmd_R45_ne295, ne295_state => state_ne295, D03_command => cmd_R45_D03, D03_state => state_D03, routeState => routes_o(44));
	route_R46 : route_45 port map(clock => clock, routeRequest => routes_i(45), ne288_command => cmd_R46_ne288, ne288_state => state_ne288, ne110_command => cmd_R46_ne110, ne110_state => state_ne110, D03_command => cmd_R46_D03, D03_state => state_D03, routeState => routes_o(45));
	route_R47 : route_46 port map(clock => clock, routeRequest => routes_i(46), ne295_command => cmd_R47_ne295, ne295_state => state_ne295, ne297_command => cmd_R47_ne297, ne297_state => state_ne297, D04_command => cmd_R47_D04, D04_state => state_D04, routeState => routes_o(46));
	route_R48 : route_47 port map(clock => clock, routeRequest => routes_i(47), ne384_command => cmd_R48_ne384, ne384_state => state_ne384, ne104_command => cmd_R48_ne104, ne104_state => state_ne104, routeState => routes_o(47));
	route_R49 : route_48 port map(clock => clock, routeRequest => routes_i(48), ne991_command => cmd_R49_ne991, ne991_state => state_ne991, ne288_command => cmd_R49_ne288, ne288_state => state_ne288, ne384_command => cmd_R49_ne384, ne384_state => state_ne384, ne110_command => cmd_R49_ne110, ne110_state => state_ne110, D01_command => cmd_R49_D01, D01_state => state_D01, D03_command => cmd_R49_D03, D03_state => state_D03, routeState => routes_o(48));
	route_R50 : route_49 port map(clock => clock, routeRequest => routes_i(49), ne295_command => cmd_R50_ne295, ne295_state => state_ne295, ne297_command => cmd_R50_ne297, ne297_state => state_ne297, D04_command => cmd_R50_D04, D04_state => state_D04, routeState => routes_o(49));
	route_R51 : route_50 port map(clock => clock, routeRequest => routes_i(50), ne297_command => cmd_R51_ne297, ne297_state => state_ne297, ne384_command => cmd_R51_ne384, ne384_state => state_ne384, D04_command => cmd_R51_D04, D04_state => state_D04, routeState => routes_o(50));
	route_R52 : route_51 port map(clock => clock, routeRequest => routes_i(51), ne400_command => cmd_R52_ne400, ne400_state => state_ne400, ne404_command => cmd_R52_ne404, ne404_state => state_ne404, D07_command => cmd_R52_D07, D07_state => state_D07, routeState => routes_o(51));
	route_R53 : route_52 port map(clock => clock, routeRequest => routes_i(52), ne400_command => cmd_R53_ne400, ne400_state => state_ne400, ne404_command => cmd_R53_ne404, ne404_state => state_ne404, D07_command => cmd_R53_D07, D07_state => state_D07, routeState => routes_o(52));
	route_R54 : route_53 port map(clock => clock, routeRequest => routes_i(53), ne400_command => cmd_R54_ne400, ne400_state => state_ne400, ne407_command => cmd_R54_ne407, ne407_state => state_ne407, D07_command => cmd_R54_D07, D07_state => state_D07, routeState => routes_o(53));
	route_R55 : route_54 port map(clock => clock, routeRequest => routes_i(54), ne61_command => cmd_R55_ne61, ne61_state => state_ne61, ne404_command => cmd_R55_ne404, ne404_state => state_ne404, ne98_command => cmd_R55_ne98, ne98_state => state_ne98, ne99_command => cmd_R55_ne99, ne99_state => state_ne99, D05_command => cmd_R55_D05, D05_state => state_D05, D08_command => cmd_R55_D08, D08_state => state_D08, routeState => routes_o(54));
	route_R56 : route_55 port map(clock => clock, routeRequest => routes_i(55), ne400_command => cmd_R56_ne400, ne400_state => state_ne400, ne407_command => cmd_R56_ne407, ne407_state => state_ne407, ne123_command => cmd_R56_ne123, ne123_state => state_ne123, D07_command => cmd_R56_D07, D07_state => state_D07, D16_command => cmd_R56_D16, D16_state => state_D16, routeState => routes_o(55));
	route_R57 : route_56 port map(clock => clock, routeRequest => routes_i(56), ne61_command => cmd_R57_ne61, ne61_state => state_ne61, ne404_command => cmd_R57_ne404, ne404_state => state_ne404, D08_command => cmd_R57_D08, D08_state => state_D08, routeState => routes_o(56));
	route_R58 : route_57 port map(clock => clock, routeRequest => routes_i(57), ne61_command => cmd_R58_ne61, ne61_state => state_ne61, ne123_command => cmd_R58_ne123, ne123_state => state_ne123, D08_command => cmd_R58_D08, D08_state => state_D08, routeState => routes_o(57));
	route_R59 : route_58 port map(clock => clock, routeRequest => routes_i(58), ne910_command => cmd_R59_ne910, ne910_state => state_ne910, ne101_command => cmd_R59_ne101, ne101_state => state_ne101, ne130_command => cmd_R59_ne130, ne130_state => state_ne130, D09_command => cmd_R59_D09, D09_state => state_D09, D10_command => cmd_R59_D10, D10_state => state_D10, routeState => routes_o(58));
	route_R60 : route_59 port map(clock => clock, routeRequest => routes_i(59), ne127_command => cmd_R60_ne127, ne127_state => state_ne127, ne135_command => cmd_R60_ne135, ne135_state => state_ne135, D24_command => cmd_R60_D24, D24_state => state_D24, routeState => routes_o(59));
	route_R61 : route_60 port map(clock => clock, routeRequest => routes_i(60), ne910_command => cmd_R61_ne910, ne910_state => state_ne910, ne130_command => cmd_R61_ne130, ne130_state => state_ne130, D10_command => cmd_R61_D10, D10_state => state_D10, routeState => routes_o(60));
	route_R62 : route_61 port map(clock => clock, routeRequest => routes_i(61), ne910_command => cmd_R62_ne910, ne910_state => state_ne910, ne135_command => cmd_R62_ne135, ne135_state => state_ne135, D10_command => cmd_R62_D10, D10_state => state_D10, routeState => routes_o(61));
	route_R63 : route_62 port map(clock => clock, routeRequest => routes_i(62), ne400_command => cmd_R63_ne400, ne400_state => state_ne400, ne993_command => cmd_R63_ne993, ne993_state => state_ne993, Sw02_command => cmd_R63_Sw02, Sw02_state => state_Sw02, routeState => routes_o(62));
	route_R64 : route_63 port map(clock => clock, routeRequest => routes_i(63), ne400_command => cmd_R64_ne400, ne400_state => state_ne400, ne993_command => cmd_R64_ne993, ne993_state => state_ne993, Sw02_command => cmd_R64_Sw02, Sw02_state => state_Sw02, routeState => routes_o(63));
	route_R65 : route_64 port map(clock => clock, routeRequest => routes_i(64), ne400_command => cmd_R65_ne400, ne400_state => state_ne400, ne992_command => cmd_R65_ne992, ne992_state => state_ne992, ne994_command => cmd_R65_ne994, ne994_state => state_ne994, Sw02_command => cmd_R65_Sw02, Sw02_state => state_Sw02, Sw01_command => cmd_R65_Sw01, Sw01_state => state_Sw01, routeState => routes_o(64));
	route_R66 : route_65 port map(clock => clock, routeRequest => routes_i(65), ne290_command => cmd_R66_ne290, ne290_state => state_ne290, ne292_command => cmd_R66_ne292, ne292_state => state_ne292, D14_command => cmd_R66_D14, D14_state => state_D14, routeState => routes_o(65));
	route_R67 : route_66 port map(clock => clock, routeRequest => routes_i(66), ne290_command => cmd_R67_ne290, ne290_state => state_ne290, ne377_command => cmd_R67_ne377, ne377_state => state_ne377, ne111_command => cmd_R67_ne111, ne111_state => state_ne111, D14_command => cmd_R67_D14, D14_state => state_D14, D15_command => cmd_R67_D15, D15_state => state_D15, routeState => routes_o(66));
	route_R68 : route_67 port map(clock => clock, routeRequest => routes_i(67), ne407_command => cmd_R68_ne407, ne407_state => state_ne407, ne122_command => cmd_R68_ne122, ne122_state => state_ne122, D16_command => cmd_R68_D16, D16_state => state_D16, routeState => routes_o(67));
	route_R69 : route_68 port map(clock => clock, routeRequest => routes_i(68), ne61_command => cmd_R69_ne61, ne61_state => state_ne61, ne407_command => cmd_R69_ne407, ne407_state => state_ne407, ne98_command => cmd_R69_ne98, ne98_state => state_ne98, ne99_command => cmd_R69_ne99, ne99_state => state_ne99, ne123_command => cmd_R69_ne123, ne123_state => state_ne123, D05_command => cmd_R69_D05, D05_state => state_D05, D08_command => cmd_R69_D08, D08_state => state_D08, D16_command => cmd_R69_D16, D16_state => state_D16, routeState => routes_o(68));
	route_R70 : route_69 port map(clock => clock, routeRequest => routes_i(69), ne63_command => cmd_R70_ne63, ne63_state => state_ne63, ne65_command => cmd_R70_ne65, ne65_state => state_ne65, D18_command => cmd_R70_D18, D18_state => state_D18, routeState => routes_o(69));
	route_R71 : route_70 port map(clock => clock, routeRequest => routes_i(70), ne63_command => cmd_R71_ne63, ne63_state => state_ne63, ne65_command => cmd_R71_ne65, ne65_state => state_ne65, D18_command => cmd_R71_D18, D18_state => state_D18, routeState => routes_o(70));
	route_R72 : route_71 port map(clock => clock, routeRequest => routes_i(71), ne63_command => cmd_R72_ne63, ne63_state => state_ne63, ne421_command => cmd_R72_ne421, ne421_state => state_ne421, ne124_command => cmd_R72_ne124, ne124_state => state_ne124, D18_command => cmd_R72_D18, D18_state => state_D18, D19_command => cmd_R72_D19, D19_state => state_D19, routeState => routes_o(71));
	route_R73 : route_72 port map(clock => clock, routeRequest => routes_i(72), ne114_command => cmd_R73_ne114, ne114_state => state_ne114, ne132_command => cmd_R73_ne132, ne132_state => state_ne132, D23_command => cmd_R73_D23, D23_state => state_D23, routeState => routes_o(72));
	route_R74 : route_73 port map(clock => clock, routeRequest => routes_i(73), ne114_command => cmd_R74_ne114, ne114_state => state_ne114, ne127_command => cmd_R74_ne127, ne127_state => state_ne127, ne129_command => cmd_R74_ne129, ne129_state => state_ne129, D23_command => cmd_R74_D23, D23_state => state_D23, D12__command => cmd_R74_D12_, D12__state => state_D12_, routeState => routes_o(73));
	route_R75 : route_74 port map(clock => clock, routeRequest => routes_i(74), ne114_command => cmd_R75_ne114, ne114_state => state_ne114, ne129_command => cmd_R75_ne129, ne129_state => state_ne129, ne130_command => cmd_R75_ne130, ne130_state => state_ne130, D23_command => cmd_R75_D23, D23_state => state_D23, D12__command => cmd_R75_D12_, D12__state => state_D12_, routeState => routes_o(74));
	route_R76 : route_75 port map(clock => clock, routeRequest => routes_i(75), ne114_command => cmd_R76_ne114, ne114_state => state_ne114, ne127_command => cmd_R76_ne127, ne127_state => state_ne127, ne129_command => cmd_R76_ne129, ne129_state => state_ne129, D23_command => cmd_R76_D23, D23_state => state_D23, D12__command => cmd_R76_D12_, D12__state => state_D12_, routeState => routes_o(75));
	route_R77 : route_76 port map(clock => clock, routeRequest => routes_i(76), ne450_command => cmd_R77_ne450, ne450_state => state_ne450, ne127_command => cmd_R77_ne127, ne127_state => state_ne127, D12__command => cmd_R77_D12_, D12__state => state_D12_, routeState => routes_o(76));
	route_R78 : route_77 port map(clock => clock, routeRequest => routes_i(77), ne114_command => cmd_R78_ne114, ne114_state => state_ne114, ne129_command => cmd_R78_ne129, ne129_state => state_ne129, ne130_command => cmd_R78_ne130, ne130_state => state_ne130, D23_command => cmd_R78_D23, D23_state => state_D23, D12__command => cmd_R78_D12_, D12__state => state_D12_, routeState => routes_o(77));
	route_R79 : route_78 port map(clock => clock, routeRequest => routes_i(78), ne450_command => cmd_R79_ne450, ne450_state => state_ne450, ne130_command => cmd_R79_ne130, ne130_state => state_ne130, D12__command => cmd_R79_D12_, D12__state => state_D12_, routeState => routes_o(78));
	route_R80 : route_79 port map(clock => clock, routeRequest => routes_i(79), ne912_command => cmd_R80_ne912, ne912_state => state_ne912, ne465_command => cmd_R80_ne465, ne465_state => state_ne465, ne131_command => cmd_R80_ne131, ne131_state => state_ne131, D20_command => cmd_R80_D20, D20_state => state_D20, D21_command => cmd_R80_D21, D21_state => state_D21, routeState => routes_o(79));
	route_R81 : route_80 port map(clock => clock, routeRequest => routes_i(80), ne912_command => cmd_R81_ne912, ne912_state => state_ne912, ne132_command => cmd_R81_ne132, ne132_state => state_ne132, D20_command => cmd_R81_D20, D20_state => state_D20, routeState => routes_o(80));
	route_R82 : route_81 port map(clock => clock, routeRequest => routes_i(81), ne910_command => cmd_R82_ne910, ne910_state => state_ne910, ne101_command => cmd_R82_ne101, ne101_state => state_ne101, ne127_command => cmd_R82_ne127, ne127_state => state_ne127, ne135_command => cmd_R82_ne135, ne135_state => state_ne135, D09_command => cmd_R82_D09, D09_state => state_D09, D10_command => cmd_R82_D10, D10_state => state_D10, D24_command => cmd_R82_D24, D24_state => state_D24, routeState => routes_o(81));
	route_R83 : route_82 port map(clock => clock, routeRequest => routes_i(82), ne127_command => cmd_R83_ne127, ne127_state => state_ne127, ne134_command => cmd_R83_ne134, ne134_state => state_ne134, D24_command => cmd_R83_D24, D24_state => state_D24, routeState => routes_o(82));
	route_R84 : route_83 port map(clock => clock, routeRequest => routes_i(83), ne65_command => cmd_R84_ne65, ne65_state => state_ne65, ne992_command => cmd_R84_ne992, ne992_state => state_ne992, Sw01_command => cmd_R84_Sw01, Sw01_state => state_Sw01, routeState => routes_o(83));
	route_R85 : route_84 port map(clock => clock, routeRequest => routes_i(84), ne65_command => cmd_R85_ne65, ne65_state => state_ne65, ne992_command => cmd_R85_ne992, ne992_state => state_ne992, Sw01_command => cmd_R85_Sw01, Sw01_state => state_Sw01, routeState => routes_o(84));
	route_R86 : route_85 port map(clock => clock, routeRequest => routes_i(85), ne400_command => cmd_R86_ne400, ne400_state => state_ne400, ne992_command => cmd_R86_ne992, ne992_state => state_ne992, ne994_command => cmd_R86_ne994, ne994_state => state_ne994, Sw02_command => cmd_R86_Sw02, Sw02_state => state_Sw02, Sw01_command => cmd_R86_Sw01, Sw01_state => state_Sw01, routeState => routes_o(85));
	route_R87 : route_86 port map(clock => clock, routeRequest => routes_i(86), ne297_command => cmd_R87_ne297, ne297_state => state_ne297, ne995_command => cmd_R87_ne995, ne995_state => state_ne995, Sw03_command => cmd_R87_Sw03, Sw03_state => state_Sw03, routeState => routes_o(86));
	route_R88 : route_87 port map(clock => clock, routeRequest => routes_i(87), ne297_command => cmd_R88_ne297, ne297_state => state_ne297, ne995_command => cmd_R88_ne995, ne995_state => state_ne995, Sw03_command => cmd_R88_Sw03, Sw03_state => state_Sw03, routeState => routes_o(87));
	route_R89 : route_88 port map(clock => clock, routeRequest => routes_i(88), ne297_command => cmd_R89_ne297, ne297_state => state_ne297, ne996_command => cmd_R89_ne996, ne996_state => state_ne996, ne997_command => cmd_R89_ne997, ne997_state => state_ne997, Sw03_command => cmd_R89_Sw03, Sw03_state => state_Sw03, Sw04_command => cmd_R89_Sw04, Sw04_state => state_Sw04, routeState => routes_o(88));
	route_R90 : route_89 port map(clock => clock, routeRequest => routes_i(89), ne292_command => cmd_R90_ne292, ne292_state => state_ne292, ne996_command => cmd_R90_ne996, ne996_state => state_ne996, Sw04_command => cmd_R90_Sw04, Sw04_state => state_Sw04, routeState => routes_o(89));
	route_R91 : route_90 port map(clock => clock, routeRequest => routes_i(90), ne297_command => cmd_R91_ne297, ne297_state => state_ne297, ne996_command => cmd_R91_ne996, ne996_state => state_ne996, ne997_command => cmd_R91_ne997, ne997_state => state_ne997, Sw03_command => cmd_R91_Sw03, Sw03_state => state_Sw03, Sw04_command => cmd_R91_Sw04, Sw04_state => state_Sw04, routeState => routes_o(90));
end Behavioral;