--  splitter.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity splitter is
		generic(
			N : natural := 316;
			N_SIGNALS : natural := 77;
			N_LEVELCROSSINGS : natural := 2;
			N_SINGLESWITCHES : natural := 22;
			N_DOUBLEWITCHES : natural := 1;
			N_ROUTES : natural := 89;
			N_TRACKCIRCUITS : natural := 47
		);
		port(
			clock : in std_logic;
			packet :  in std_logic_vector(N-1 downto 0);
			processing :  in std_logic;
			processed :  out std_logic;
			ocupation :  out std_logic_vector(N_TRACKCIRCUITS-1 downto 0);
			signals :  out signals_type;
			routes : out std_logic_vector(N_ROUTES-1 downto 0);
			levelCrossings : out std_logic_vector(N_LEVELCROSSINGS-1 downto 0);
			singleSwitches : out std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			doubleSwitches : out dSwitch_type;
			reset : in std_logic
		);
	end entity splitter;
architecture Behavioral of splitter is
	Signal tc_s : std_logic_vector(47-1 downto 0);
	Signal sig_s_i,sig_s_o : signals_type;
	Signal rt_s_i,rt_s_o : std_logic_vector(89-1 downto 0);
	Signal lc_s_i,lc_s_o : std_logic_vector(2-1 downto 0);
	Signal ssw_s_i,ssw_s_o : std_logic_vector(22-1 downto 0);
	Signal dsw_s_i,dsw_s_o : dSwitch_type;
begin
	process(clock,reset)
	begin
		if (clock = '1' and clock'Event) then
			if (reset = '1') then
				ocupation <= "00000000000000000000000000000000000000000000000";
				signals.lsb <= "00000000000000000000000000000000000000000000000000000000000000000000000000000";
				signals.msb <= "00000000000000000000000000000000000000000000000000000000000000000000000000000";
				routes <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
				levelCrossings <= "00";
				singleSwitches <= "0000000000000000000000";
				doubleSwitches.lsb <= '0';
				doubleSwitches.msb <= '0';
				processed <= '0';
			else
				processed <= processing;
				if processing = '1' then
					ocupation(0) <= packet(315);
					ocupation(1) <= packet(314);
					ocupation(2) <= packet(313);
					ocupation(3) <= packet(312);
					ocupation(4) <= packet(311);
					ocupation(5) <= packet(310);
					ocupation(6) <= packet(309);
					ocupation(7) <= packet(308);
					ocupation(8) <= packet(307);
					ocupation(9) <= packet(306);
					ocupation(10) <= packet(305);
					ocupation(11) <= packet(304);
					ocupation(12) <= packet(303);
					ocupation(13) <= packet(302);
					ocupation(14) <= packet(301);
					ocupation(15) <= packet(300);
					ocupation(16) <= packet(299);
					ocupation(17) <= packet(298);
					ocupation(18) <= packet(297);
					ocupation(19) <= packet(296);
					ocupation(20) <= packet(295);
					ocupation(21) <= packet(294);
					ocupation(22) <= packet(293);
					ocupation(23) <= packet(292);
					ocupation(24) <= packet(291);
					ocupation(25) <= packet(290);
					ocupation(26) <= packet(289);
					ocupation(27) <= packet(288);
					ocupation(28) <= packet(287);
					ocupation(29) <= packet(286);
					ocupation(30) <= packet(285);
					ocupation(31) <= packet(284);
					ocupation(32) <= packet(283);
					ocupation(33) <= packet(282);
					ocupation(34) <= packet(281);
					ocupation(35) <= packet(280);
					ocupation(36) <= packet(279);
					ocupation(37) <= packet(278);
					ocupation(38) <= packet(277);
					ocupation(39) <= packet(276);
					ocupation(40) <= packet(275);
					ocupation(41) <= packet(274);
					ocupation(42) <= packet(273);
					ocupation(43) <= packet(272);
					ocupation(44) <= packet(271);
					ocupation(45) <= packet(270);
					ocupation(46) <= packet(269);
					routes(0) <= packet(268);
					routes(1) <= packet(267);
					routes(2) <= packet(266);
					routes(3) <= packet(265);
					routes(4) <= packet(264);
					routes(5) <= packet(263);
					routes(6) <= packet(262);
					routes(7) <= packet(261);
					routes(8) <= packet(260);
					routes(9) <= packet(259);
					routes(10) <= packet(258);
					routes(11) <= packet(257);
					routes(12) <= packet(256);
					routes(13) <= packet(255);
					routes(14) <= packet(254);
					routes(15) <= packet(253);
					routes(16) <= packet(252);
					routes(17) <= packet(251);
					routes(18) <= packet(250);
					routes(19) <= packet(249);
					routes(20) <= packet(248);
					routes(21) <= packet(247);
					routes(22) <= packet(246);
					routes(23) <= packet(245);
					routes(24) <= packet(244);
					routes(25) <= packet(243);
					routes(26) <= packet(242);
					routes(27) <= packet(241);
					routes(28) <= packet(240);
					routes(29) <= packet(239);
					routes(30) <= packet(238);
					routes(31) <= packet(237);
					routes(32) <= packet(236);
					routes(33) <= packet(235);
					routes(34) <= packet(234);
					routes(35) <= packet(233);
					routes(36) <= packet(232);
					routes(37) <= packet(231);
					routes(38) <= packet(230);
					routes(39) <= packet(229);
					routes(40) <= packet(228);
					routes(41) <= packet(227);
					routes(42) <= packet(226);
					routes(43) <= packet(225);
					routes(44) <= packet(224);
					routes(45) <= packet(223);
					routes(46) <= packet(222);
					routes(47) <= packet(221);
					routes(48) <= packet(220);
					routes(49) <= packet(219);
					routes(50) <= packet(218);
					routes(51) <= packet(217);
					routes(52) <= packet(216);
					routes(53) <= packet(215);
					routes(54) <= packet(214);
					routes(55) <= packet(213);
					routes(56) <= packet(212);
					routes(57) <= packet(211);
					routes(58) <= packet(210);
					routes(59) <= packet(209);
					routes(60) <= packet(208);
					routes(61) <= packet(207);
					routes(62) <= packet(206);
					routes(63) <= packet(205);
					routes(64) <= packet(204);
					routes(65) <= packet(203);
					routes(66) <= packet(202);
					routes(67) <= packet(201);
					routes(68) <= packet(200);
					routes(69) <= packet(199);
					routes(70) <= packet(198);
					routes(71) <= packet(197);
					routes(72) <= packet(196);
					routes(73) <= packet(195);
					routes(74) <= packet(194);
					routes(75) <= packet(193);
					routes(76) <= packet(192);
					routes(77) <= packet(191);
					routes(78) <= packet(190);
					routes(79) <= packet(189);
					routes(80) <= packet(188);
					routes(81) <= packet(187);
					routes(82) <= packet(186);
					routes(83) <= packet(185);
					routes(84) <= packet(184);
					routes(85) <= packet(183);
					routes(86) <= packet(182);
					routes(87) <= packet(181);
					routes(88) <= packet(180);
					signals.msb(0) <= packet(179);
					signals.lsb(0) <= packet(178);
					signals.msb(1) <= packet(177);
					signals.lsb(1) <= packet(176);
					signals.msb(2) <= packet(175);
					signals.lsb(2) <= packet(174);
					signals.msb(3) <= packet(173);
					signals.lsb(3) <= packet(172);
					signals.msb(4) <= packet(171);
					signals.lsb(4) <= packet(170);
					signals.msb(5) <= packet(169);
					signals.lsb(5) <= packet(168);
					signals.msb(6) <= packet(167);
					signals.lsb(6) <= packet(166);
					signals.msb(7) <= packet(165);
					signals.lsb(7) <= packet(164);
					signals.msb(8) <= packet(163);
					signals.lsb(8) <= packet(162);
					signals.msb(9) <= packet(161);
					signals.lsb(9) <= packet(160);
					signals.msb(10) <= packet(159);
					signals.lsb(10) <= packet(158);
					signals.msb(11) <= packet(157);
					signals.lsb(11) <= packet(156);
					signals.msb(12) <= packet(155);
					signals.lsb(12) <= packet(154);
					signals.msb(13) <= packet(153);
					signals.lsb(13) <= packet(152);
					signals.msb(14) <= packet(151);
					signals.lsb(14) <= packet(150);
					signals.msb(15) <= packet(149);
					signals.lsb(15) <= packet(148);
					signals.msb(16) <= packet(147);
					signals.lsb(16) <= packet(146);
					signals.msb(17) <= packet(145);
					signals.lsb(17) <= packet(144);
					signals.msb(18) <= packet(143);
					signals.lsb(18) <= packet(142);
					signals.msb(19) <= packet(141);
					signals.lsb(19) <= packet(140);
					signals.msb(20) <= packet(139);
					signals.lsb(20) <= packet(138);
					signals.msb(21) <= packet(137);
					signals.lsb(21) <= packet(136);
					signals.msb(22) <= packet(135);
					signals.lsb(22) <= packet(134);
					signals.msb(23) <= packet(133);
					signals.lsb(23) <= packet(132);
					signals.msb(24) <= packet(131);
					signals.lsb(24) <= packet(130);
					signals.msb(25) <= packet(129);
					signals.lsb(25) <= packet(128);
					signals.msb(26) <= packet(127);
					signals.lsb(26) <= packet(126);
					signals.msb(27) <= packet(125);
					signals.lsb(27) <= packet(124);
					signals.msb(28) <= packet(123);
					signals.lsb(28) <= packet(122);
					signals.msb(29) <= packet(121);
					signals.lsb(29) <= packet(120);
					signals.msb(30) <= packet(119);
					signals.lsb(30) <= packet(118);
					signals.msb(31) <= packet(117);
					signals.lsb(31) <= packet(116);
					signals.msb(32) <= packet(115);
					signals.lsb(32) <= packet(114);
					signals.msb(33) <= packet(113);
					signals.lsb(33) <= packet(112);
					signals.msb(34) <= packet(111);
					signals.lsb(34) <= packet(110);
					signals.msb(35) <= packet(109);
					signals.lsb(35) <= packet(108);
					signals.msb(36) <= packet(107);
					signals.lsb(36) <= packet(106);
					signals.msb(37) <= packet(105);
					signals.lsb(37) <= packet(104);
					signals.msb(38) <= packet(103);
					signals.lsb(38) <= packet(102);
					signals.msb(39) <= packet(101);
					signals.lsb(39) <= packet(100);
					signals.msb(40) <= packet(99);
					signals.lsb(40) <= packet(98);
					signals.msb(41) <= packet(97);
					signals.lsb(41) <= packet(96);
					signals.msb(42) <= packet(95);
					signals.lsb(42) <= packet(94);
					signals.msb(43) <= packet(93);
					signals.lsb(43) <= packet(92);
					signals.msb(44) <= packet(91);
					signals.lsb(44) <= packet(90);
					signals.msb(45) <= packet(89);
					signals.lsb(45) <= packet(88);
					signals.msb(46) <= packet(87);
					signals.lsb(46) <= packet(86);
					signals.msb(47) <= packet(85);
					signals.lsb(47) <= packet(84);
					signals.msb(48) <= packet(83);
					signals.lsb(48) <= packet(82);
					signals.msb(49) <= packet(81);
					signals.lsb(49) <= packet(80);
					signals.msb(50) <= packet(79);
					signals.lsb(50) <= packet(78);
					signals.msb(51) <= packet(77);
					signals.lsb(51) <= packet(76);
					signals.msb(52) <= packet(75);
					signals.lsb(52) <= packet(74);
					signals.msb(53) <= packet(73);
					signals.lsb(53) <= packet(72);
					signals.msb(54) <= packet(71);
					signals.lsb(54) <= packet(70);
					signals.msb(55) <= packet(69);
					signals.lsb(55) <= packet(68);
					signals.msb(56) <= packet(67);
					signals.lsb(56) <= packet(66);
					signals.msb(57) <= packet(65);
					signals.lsb(57) <= packet(64);
					signals.msb(58) <= packet(63);
					signals.lsb(58) <= packet(62);
					signals.msb(59) <= packet(61);
					signals.lsb(59) <= packet(60);
					signals.msb(60) <= packet(59);
					signals.lsb(60) <= packet(58);
					signals.msb(61) <= packet(57);
					signals.lsb(61) <= packet(56);
					signals.msb(62) <= packet(55);
					signals.lsb(62) <= packet(54);
					signals.msb(63) <= packet(53);
					signals.lsb(63) <= packet(52);
					signals.msb(64) <= packet(51);
					signals.lsb(64) <= packet(50);
					signals.msb(65) <= packet(49);
					signals.lsb(65) <= packet(48);
					signals.msb(66) <= packet(47);
					signals.lsb(66) <= packet(46);
					signals.msb(67) <= packet(45);
					signals.lsb(67) <= packet(44);
					signals.msb(68) <= packet(43);
					signals.lsb(68) <= packet(42);
					signals.msb(69) <= packet(41);
					signals.lsb(69) <= packet(40);
					signals.msb(70) <= packet(39);
					signals.lsb(70) <= packet(38);
					signals.msb(71) <= packet(37);
					signals.lsb(71) <= packet(36);
					signals.msb(72) <= packet(35);
					signals.lsb(72) <= packet(34);
					signals.msb(73) <= packet(33);
					signals.lsb(73) <= packet(32);
					signals.msb(74) <= packet(31);
					signals.lsb(74) <= packet(30);
					signals.msb(75) <= packet(29);
					signals.lsb(75) <= packet(28);
					signals.msb(76) <= packet(27);
					signals.lsb(76) <= packet(26);
					levelCrossings(0) <= packet(25);
					levelCrossings(1) <= packet(24);
					singleSwitches(0) <= packet(23);
					singleSwitches(1) <= packet(22);
					singleSwitches(2) <= packet(21);
					singleSwitches(3) <= packet(20);
					singleSwitches(4) <= packet(19);
					singleSwitches(5) <= packet(18);
					singleSwitches(6) <= packet(17);
					singleSwitches(7) <= packet(16);
					singleSwitches(8) <= packet(15);
					singleSwitches(9) <= packet(14);
					singleSwitches(10) <= packet(13);
					singleSwitches(11) <= packet(12);
					singleSwitches(12) <= packet(11);
					singleSwitches(13) <= packet(10);
					singleSwitches(14) <= packet(9);
					singleSwitches(15) <= packet(8);
					singleSwitches(16) <= packet(7);
					singleSwitches(17) <= packet(6);
					singleSwitches(18) <= packet(5);
					singleSwitches(19) <= packet(4);
					singleSwitches(20) <= packet(3);
					singleSwitches(21) <= packet(2);
					doubleSwitches.lsb <= packet(1);
					doubleSwitches.msb <= packet(0);
				end if;
			end if;
		end if;
	end process;
end Behavioral;