--  railwaySignal_43.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
--Declare the package
use work.my_package.all;
	entity railwaySignal_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R33_command : in routeCommands;
			R25_command : in routeCommands;
			Lc04_state : in hex_char;
			--Ocupation level 0
			track_ne100 : in hex_char;
			correspondence_X53 : out hex_char;
			--Ocupation level 1
			track_ne992 : in hex_char;
			correspondence_S120 : in hex_char;
			--Ocupation level 2
			track_ne994 : in hex_char;
			track_ne65 : in hex_char;
			track_ne400 : in hex_char;
			correspondence_C94 : in hex_char;
			correspondence_S74 : in hex_char;
			Sw01_state : in hex_char;
			Sw05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end entity railwaySignal_43;
architecture Behavioral of railwaySignal_43 is
	component flipFlop is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			Q : out std_logic := '0'
		);
	end component flipFlop;
	signal restart : std_logic := '1';
	signal Q : std_logic_vector(30 downto 0) := (others => '0');
	signal clock_in : std_logic_vector(30 downto 0) := (others => '0');
	signal timeout : std_logic := '0';
	signal commandState : routeCommands := RELEASE;
	signal lockStateIn : objectLock := RELEASED;
	signal lockStateOut : objectLock := RELEASED;
	signal aspectStateIn : signalStates := RED;
	signal aspectStateOut : signalStates := RED;
	signal correspondenceState : signalStates := RED;
	signal path : integer := 0;
	signal Lc04_position : levelCrossingStates := UP;
	signal Lc04_lock : objectLock := RELEASED;
	--Ocupation level 1
	signal ne992_state : nodeStates := FREE;
	signal ne992_lock : objectLock := RELEASED;
	signal S120_aspect : signalStates;
	signal S120_lock : objectLock := RELEASED;
	--Ocupation level 2
	signal ne994_state : nodeStates := FREE;
	signal ne994_lock : objectLock := RELEASED;
	signal ne65_state : nodeStates := FREE;
	signal ne65_lock : objectLock := RELEASED;
	signal ne400_state : nodeStates := FREE;
	signal ne400_lock : objectLock := RELEASED;
	signal C94_aspect : signalStates;
	signal C94_lock : objectLock := RELEASED;
	signal S74_aspect : signalStates;
	signal S74_lock : objectLock := RELEASED;
	signal Sw01_position : singleSwitchStates := NORMAL;
	signal Sw05_position : singleSwitchStates := NORMAL;
	signal Sw01_lock : objectLock := RELEASED;
	signal Sw05_lock : objectLock := RELEASED;
begin
	clock_in(0) <= clock;
	lockStateIn <= objectLock'val(to_integer(unsigned(hex_to_slv(indication)(0 to 1))));
	aspectStateIn <= signalStates'val(to_integer(unsigned(hex_to_slv(indication)(2 to 3))));
	command <= slv_to_hex(std_logic_vector(to_unsigned(objectLock'pos(lockStateOut), 2) & to_unsigned(signalStates'pos(aspectStateOut), 2)));
	correspondence_X53 <= slv_to_hex(std_logic_vector(to_unsigned(objectLock'pos(lockStateOut), 2) & to_unsigned(signalStates'pos(correspondenceState), 2)));
	Lc04_position <= levelCrossingStates'val(to_integer(unsigned(hex_to_slv(Lc04_state)(2 to 3))));
	Lc04_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(Lc04_state)(0 to 1))));
	--Ocupation level 1
	ne992_state <= nodeStates'val(to_integer(unsigned(hex_to_slv(track_ne992)(2 to 3))));
	ne992_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(track_ne992)(0 to 1))));
	S120_aspect <= signalStates'val(to_integer(unsigned(hex_to_slv(correspondence_S120)(2 to 3))));
	S120_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(correspondence_S120)(0 to 1))));
	--Ocupation level 2
	ne994_state <= nodeStates'val(to_integer(unsigned(hex_to_slv(track_ne994)(2 to 3))));
	ne994_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(track_ne994)(0 to 1))));
	ne65_state <= nodeStates'val(to_integer(unsigned(hex_to_slv(track_ne65)(2 to 3))));
	ne65_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(track_ne65)(0 to 1))));
	ne400_state <= nodeStates'val(to_integer(unsigned(hex_to_slv(track_ne400)(2 to 3))));
	ne400_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(track_ne400)(0 to 1))));
	C94_aspect <= signalStates'val(to_integer(unsigned(hex_to_slv(correspondence_C94)(2 to 3))));
	C94_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(correspondence_C94)(0 to 1))));
	S74_aspect <= signalStates'val(to_integer(unsigned(hex_to_slv(correspondence_S74)(2 to 3))));
	S74_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(correspondence_S74)(0 to 1))));
	Sw01_position <= singleSwitchStates'val(to_integer(unsigned(hex_to_slv(Sw01_state)(2 to 3))));
	Sw05_position <= singleSwitchStates'val(to_integer(unsigned(hex_to_slv(Sw05_state)(2 to 3))));
	Sw01_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(Sw01_state)(0 to 1))));
	Sw05_lock <= objectLock'val(to_integer(unsigned(hex_to_slv(Sw05_state)(0 to 1))));
	gen : for i in 0 to 29 generate
		inst: flipFlop port map(Q(i),restart,Q(i+1));
	end generate;

	process(timeout,R33_command,R25_command)
	begin
		if (timeout = '1') then
			commandState <= RELEASE;
		else
			if (R33_command = RELEASE and R25_command = RELEASE) then
				commandState <= RELEASE;
			end if;
			if (R33_command = RESERVE or R25_command = RESERVE) then
				commandState <= RESERVE;
			end if;
			if (R33_command = LOCK or R25_command = LOCK) then
				commandState <= LOCK;
			end if;
		end if;
	end process;

	process(commandState)
	begin
		case commandState is
			when RELEASE => -- AUTOMATIC
				lockStateOut <= RELEASED;
			when RESERVE => -- DONT CHANGE
				lockStateOut <= RESERVED;
			when LOCK => -- DONT CHANGE
				lockStateOut <= LOCKED;
			when others =>
				lockStateOut <= LOCKED;
		end case;
	end process;

	process(commandState,Sw01_position,Sw01_position,Sw05_position)
	begin
		case commandState is
			when RELEASE =>
				if ((Sw01_position = NORMAL and Sw01_position = REVERSE and Sw05_position = REVERSE and Lc04_position = DOWN) or (Sw01_position = NORMAL and Sw01_position = REVERSE and Sw05_position = REVERSE and Lc04_position = DOWN)) then
					if (Sw01_position = NORMAL and Sw01_position = REVERSE and Sw05_position = REVERSE and Lc04_position = DOWN) then
						path <= 1;
					end if;
					if (Sw01_position = NORMAL and Sw01_position = REVERSE and Sw05_position = REVERSE and Lc04_position = DOWN) then
						path <= 2;
					end if;
				else
					path <= 0;
				end if;
			when RESERVE =>
				path <= 3;
			when LOCK =>
				path <= 0;
			when others =>
				path <= 0;
		end case;
	end process;

	process(path,ne992_state,S120_aspect)
	begin
		case path is
			when 0 =>
				aspectStateOut <= RED;
			when 1 =>
				if (ne992_state = OCCUPIED or ne992_lock = LOCKED) then
					aspectStateOut <= RED;
				else
					if (S120_aspect = RED) then
						aspectStateOut <= DOUBLE_YELLOW;
					end if;
					if (S120_aspect = DOUBLE_YELLOW) then
						aspectStateOut <= YELLOW;
					end if;
					if (S120_aspect = YELLOW) then
						aspectStateOut <= GREEN;
					end if;
					if (S120_aspect = GREEN) then
						aspectStateOut <= GREEN;
					end if;
				end if;
			when 2 =>
				if (ne992_state = OCCUPIED or ne992_lock = LOCKED) then
					aspectStateOut <= RED;
				else
					if (S120_aspect = RED) then
						aspectStateOut <= DOUBLE_YELLOW;
					end if;
					if (S120_aspect = DOUBLE_YELLOW) then
						aspectStateOut <= YELLOW;
					end if;
					if (S120_aspect = YELLOW) then
						aspectStateOut <= GREEN;
					end if;
					if (S120_aspect = GREEN) then
						aspectStateOut <= GREEN;
					end if;
				end if;
			when 3 =>
				aspectStateOut <= GREEN;
			when others =>
				aspectStateOut <= RED;
		end case;
	end process;

	process(clock,reset,Q,restart)
	begin
		if (reset = '1' or Q = "010100110111001001001110000000") then
			timeout <= '1';
		end if;
		if (restart = '1') then
			timeout <= '0';
		end if;
	end process;

	process(timeout,aspectStateOut,aspectStateIn)
	begin
		if(aspectStateOut = RED and aspectStateIn = RED) then
			correspondenceState <= RED;
			restart <= '1';
		end if;
		if(aspectStateOut = GREEN and aspectStateIn = GREEN) then
			correspondenceState <= GREEN;
			restart <= '1';
		end if;
		if(aspectStateOut = DOUBLE_YELLOW and aspectStateIn = DOUBLE_YELLOW) then
			correspondenceState <= DOUBLE_YELLOW;
			restart <= '1';
		end if;
		if(aspectStateOut = YELLOW and aspectStateIn = YELLOW) then
			correspondenceState <= YELLOW;
			restart <= '1';
		end if;
	end process;
end Behavioral;