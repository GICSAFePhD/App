--  route_52.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity route_52 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne29_state : in nodeStates;
			ne29_command : out routeCommands;
			ne30_state : in nodeStates;
			ne30_command : out routeCommands;
			Sw08_state : in singleSwitchStates;
			Sw08_command : out routeCommands;
			routeState : out std_logic
		);
	end entity route_52;
architecture Behavioral of route_52 is
begin
	routeState <= '0';
end Behavioral;