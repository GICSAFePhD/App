--  network.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
--Declare the package
use work.my_package.all;
	entity network is
		generic(
			N_TRACKCIRCUITS : natural := 47;
			N_ROUTES : natural := 89;
			N_SIGNALS : natural := 77;
			N_LEVELCROSSINGS : natural := 2;
			N_SINGLESWITCHES : natural := 22;
			N_DOUBLESWITCHES : natural := 1;
			N : natural := 238
		);
		port(
			clock : in std_logic;
			processing : in std_logic;
			processed : out std_logic;
			tracks_i : in hex_array(N_TRACKCIRCUITS-1 downto 0);
			tracks_o : out hex_array(N_TRACKCIRCUITS-1 downto 0);
			signals_i : in hex_array(N_SIGNALS-1 downto 0);
			signals_o : out hex_array(N_SIGNALS-1 downto 0);
			routes_i : in hex_array(N_ROUTES-1 downto 0);
			routes_o : out hex_array(N_ROUTES-1 downto 0);
			levelCrossings_i : in hex_array(N_LEVELCROSSINGS-1 downto 0);
			levelCrossings_o : out hex_array(N_LEVELCROSSINGS-1 downto 0);
			singleSwitches_i : in hex_array(N_SINGLESWITCHES-1 downto 0);
			singleSwitches_o : out hex_array(N_SINGLESWITCHES-1 downto 0);
			doubleSwitches_i : in hex_char;
			doubleSwitches_o : out hex_char;
			reset : in std_logic
		);
	end entity network;
architecture Behavioral of network is
	component levelCrossing_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			track_ne98 : in hex_char;
			track_ne996 : in hex_char;
			track_ne99 : in hex_char;
			R30_command : in routeCommands;
			R31_command : in routeCommands;
			R34_command : in routeCommands;
			R51_command : in routeCommands;
			R64_command : in routeCommands;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component levelCrossing_0;
	component levelCrossing_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			track_ne100 : in hex_char;
			track_ne992 : in hex_char;
			track_ne101 : in hex_char;
			R32_command : in routeCommands;
			R33_command : in routeCommands;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component levelCrossing_1;
	component singleSwitch_0 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R20_command : in routeCommands := RELEASE;
			R39_command : in routeCommands := RELEASE;
			R40_command : in routeCommands := RELEASE;
			R41_command : in routeCommands := RELEASE;
			R60_command : in routeCommands := RELEASE;
			R1_command : in routeCommands := RELEASE;
			R22_command : in routeCommands := RELEASE;
			R46_command : in routeCommands := RELEASE;
			R2_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_0;
	component singleSwitch_1 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R51_command : in routeCommands := RELEASE;
			R53_command : in routeCommands := RELEASE;
			R54_command : in routeCommands := RELEASE;
			R64_command : in routeCommands := RELEASE;
			R49_command : in routeCommands := RELEASE;
			R35_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_1;
	component singleSwitch_2 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R34_command : in routeCommands := RELEASE;
			R35_command : in routeCommands := RELEASE;
			R36_command : in routeCommands := RELEASE;
			R51_command : in routeCommands := RELEASE;
			R64_command : in routeCommands := RELEASE;
			R65_command : in routeCommands := RELEASE;
			R49_command : in routeCommands := RELEASE;
			R4_command : in routeCommands := RELEASE;
			R30_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_2;
	component singleSwitch_3 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R4_command : in routeCommands := RELEASE;
			R65_command : in routeCommands := RELEASE;
			R66_command : in routeCommands := RELEASE;
			R67_command : in routeCommands := RELEASE;
			R36_command : in routeCommands := RELEASE;
			R80_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_3;
	component singleSwitch_4 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R79_command : in routeCommands := RELEASE;
			R80_command : in routeCommands := RELEASE;
			R81_command : in routeCommands := RELEASE;
			R84_command : in routeCommands := RELEASE;
			R66_command : in routeCommands := RELEASE;
			R33_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_4;
	component singleSwitch_5 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R55_command : in routeCommands := RELEASE;
			R57_command : in routeCommands := RELEASE;
			R58_command : in routeCommands := RELEASE;
			R77_command : in routeCommands := RELEASE;
			R69_command : in routeCommands := RELEASE;
			R70_command : in routeCommands := RELEASE;
			R6_command : in routeCommands := RELEASE;
			R7_command : in routeCommands := RELEASE;
			R38_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_5;
	component singleSwitch_6 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R26_command : in routeCommands := RELEASE;
			R37_command : in routeCommands := RELEASE;
			R38_command : in routeCommands := RELEASE;
			R55_command : in routeCommands := RELEASE;
			R77_command : in routeCommands := RELEASE;
			R69_command : in routeCommands := RELEASE;
			R70_command : in routeCommands := RELEASE;
			R6_command : in routeCommands := RELEASE;
			R7_command : in routeCommands := RELEASE;
			R8_command : in routeCommands := RELEASE;
			R32_command : in routeCommands := RELEASE;
			R28_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_6;
	component singleSwitch_7 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R8_command : in routeCommands := RELEASE;
			R28_command : in routeCommands := RELEASE;
			R75_command : in routeCommands := RELEASE;
			R76_command : in routeCommands := RELEASE;
			R68_command : in routeCommands := RELEASE;
			R37_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_7;
	component singleSwitch_8 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R27_command : in routeCommands := RELEASE;
			R68_command : in routeCommands := RELEASE;
			R69_command : in routeCommands := RELEASE;
			R70_command : in routeCommands := RELEASE;
			R71_command : in routeCommands := RELEASE;
			R73_command : in routeCommands := RELEASE;
			R57_command : in routeCommands := RELEASE;
			R76_command : in routeCommands := RELEASE;
			R10_command : in routeCommands := RELEASE;
			R16_command : in routeCommands := RELEASE;
			R56_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_8;
	component singleSwitch_9 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R41_command : in routeCommands := RELEASE;
			R43_command : in routeCommands := RELEASE;
			R44_command : in routeCommands := RELEASE;
			R60_command : in routeCommands := RELEASE;
			R39_command : in routeCommands := RELEASE;
			R46_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_9;
	component singleSwitch_10 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R2_command : in routeCommands := RELEASE;
			R22_command : in routeCommands := RELEASE;
			R61_command : in routeCommands := RELEASE;
			R62_command : in routeCommands := RELEASE;
			R40_command : in routeCommands := RELEASE;
			R88_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_10;
	component singleSwitch_11 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R21_command : in routeCommands := RELEASE;
			R87_command : in routeCommands := RELEASE;
			R88_command : in routeCommands := RELEASE;
			R89_command : in routeCommands := RELEASE;
			R61_command : in routeCommands := RELEASE;
			R31_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_11;
	component singleSwitch_12 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R11_command : in routeCommands := RELEASE;
			R42_command : in routeCommands := RELEASE;
			R45_command : in routeCommands := RELEASE;
			R46_command : in routeCommands := RELEASE;
			R47_command : in routeCommands := RELEASE;
			R43_command : in routeCommands := RELEASE;
			R44_command : in routeCommands := RELEASE;
			R85_command : in routeCommands := RELEASE;
			R89_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_12;
	component singleSwitch_13 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R85_command : in routeCommands := RELEASE;
			R86_command : in routeCommands := RELEASE;
			R87_command : in routeCommands := RELEASE;
			R89_command : in routeCommands := RELEASE;
			R45_command : in routeCommands := RELEASE;
			R31_command : in routeCommands := RELEASE;
			R11_command : in routeCommands := RELEASE;
			R42_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_13;
	component singleSwitch_14 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R2_command : in routeCommands := RELEASE;
			R3_command : in routeCommands := RELEASE;
			R12_command : in routeCommands := RELEASE;
			R62_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_14;
	component singleSwitch_15 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R11_command : in routeCommands := RELEASE;
			R42_command : in routeCommands := RELEASE;
			R59_command : in routeCommands := RELEASE;
			R60_command : in routeCommands := RELEASE;
			R44_command : in routeCommands := RELEASE;
			R47_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_15;
	component singleSwitch_16 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R13_command : in routeCommands := RELEASE;
			R48_command : in routeCommands := RELEASE;
			R49_command : in routeCommands := RELEASE;
			R50_command : in routeCommands := RELEASE;
			R52_command : in routeCommands := RELEASE;
			R53_command : in routeCommands := RELEASE;
			R54_command : in routeCommands := RELEASE;
			R81_command : in routeCommands := RELEASE;
			R82_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_16;
	component singleSwitch_17 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R81_command : in routeCommands := RELEASE;
			R82_command : in routeCommands := RELEASE;
			R83_command : in routeCommands := RELEASE;
			R84_command : in routeCommands := RELEASE;
			R48_command : in routeCommands := RELEASE;
			R33_command : in routeCommands := RELEASE;
			R13_command : in routeCommands := RELEASE;
			R52_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_17;
	component singleSwitch_18 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R13_command : in routeCommands := RELEASE;
			R52_command : in routeCommands := RELEASE;
			R63_command : in routeCommands := RELEASE;
			R64_command : in routeCommands := RELEASE;
			R54_command : in routeCommands := RELEASE;
			R50_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_18;
	component singleSwitch_19 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R4_command : in routeCommands := RELEASE;
			R5_command : in routeCommands := RELEASE;
			R14_command : in routeCommands := RELEASE;
			R67_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_19;
	component singleSwitch_20 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R8_command : in routeCommands := RELEASE;
			R9_command : in routeCommands := RELEASE;
			R15_command : in routeCommands := RELEASE;
			R75_command : in routeCommands := RELEASE;
			R37_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_20;
	component singleSwitch_21 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R16_command : in routeCommands := RELEASE;
			R56_command : in routeCommands := RELEASE;
			R77_command : in routeCommands := RELEASE;
			R78_command : in routeCommands := RELEASE;
			R58_command : in routeCommands := RELEASE;
			R69_command : in routeCommands := RELEASE;
			R6_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_21;
	component doubleSwitch_0 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R6_command : in routeCommands := RELEASE;
			R7_command : in routeCommands := RELEASE;
			R69_command : in routeCommands := RELEASE;
			R70_command : in routeCommands := RELEASE;
			R71_command : in routeCommands := RELEASE;
			R72_command : in routeCommands := RELEASE;
			R73_command : in routeCommands := RELEASE;
			R74_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component doubleSwitch_0;
	component railwaySignal_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R20_command : in routeCommands;
			R41_command : in routeCommands;
			R60_command : in routeCommands;
			--Ocupation level 0
			track_ne991 : in hex_char;
			correspondence_T01 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_0;
	component railwaySignal_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R1_command : in routeCommands;
			--Ocupation level 0
			track_ne991 : in hex_char;
			correspondence_T02 : out hex_char;
			correspondence_S64 : in hex_char;
			--Ocupation level 2
			track_ne290 : in hex_char;
			track_ne288 : in hex_char;
			correspondence_S69 : in hex_char;
			correspondence_S86 : in hex_char;
			D01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_1;
	component railwaySignal_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			R1_command : in routeCommands;
			--Ocupation level 0
			track_ne991 : in hex_char;
			correspondence_S64 : out hex_char;
			--Ocupation level 1
			track_ne288 : in hex_char;
			track_ne290 : in hex_char;
			correspondence_S69 : in hex_char;
			correspondence_S86 : in hex_char;
			D01_state : in hex_char;
			--Ocupation level 2
			track_ne295 : in hex_char;
			track_ne110 : in hex_char;
			track_ne292 : in hex_char;
			track_ne111 : in hex_char;
			track_ne377 : in hex_char;
			correspondence_C70 : in hex_char;
			correspondence_B68 : in hex_char;
			correspondence_J36 : in hex_char;
			correspondence_T03 : in hex_char;
			D03_state : in hex_char;
			D14_state : in hex_char;
			D15_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_2;
	component railwaySignal_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R35_command : in routeCommands;
			--Ocupation level 0
			track_ne61 : in hex_char;
			correspondence_S78 : out hex_char;
			--Ocupation level 1
			track_ne404 : in hex_char;
			track_ne123 : in hex_char;
			correspondence_C73 : in hex_char;
			correspondence_B77 : in hex_char;
			D08_state : in hex_char;
			--Ocupation level 2
			track_ne400 : in hex_char;
			track_ne407 : in hex_char;
			correspondence_S123 : in hex_char;
			D07_state : in hex_char;
			D16_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_3;
	component railwaySignal_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R34_command : in routeCommands;
			R4_command : in routeCommands;
			R65_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne63 : in hex_char;
			correspondence_C54 : out hex_char;
			--Ocupation level 1
			track_ne99 : in hex_char;
			track_ne98 : in hex_char;
			correspondence_X51 : in hex_char;
			D05_state : in hex_char;
			--Ocupation level 2
			track_ne996 : in hex_char;
			correspondence_S129 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_4;
	component railwaySignal_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R66_command : in routeCommands;
			R67_command : in routeCommands;
			R36_command : in routeCommands;
			--Ocupation level 0
			track_ne63 : in hex_char;
			correspondence_S95 : out hex_char;
			--Ocupation level 1
			track_ne65 : in hex_char;
			track_ne124 : in hex_char;
			track_ne421 : in hex_char;
			correspondence_C119 : in hex_char;
			correspondence_T05 : in hex_char;
			D18_state : in hex_char;
			D19_state : in hex_char;
			--Ocupation level 2
			track_ne992 : in hex_char;
			correspondence_J40 : in hex_char;
			Sw01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_5;
	component railwaySignal_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R65_command : in routeCommands;
			R80_command : in routeCommands;
			--Ocupation level 0
			track_ne65 : in hex_char;
			correspondence_C94 : out hex_char;
			--Ocupation level 1
			track_ne63 : in hex_char;
			correspondence_C54 : in hex_char;
			D18_state : in hex_char;
			--Ocupation level 2
			track_ne98 : in hex_char;
			track_ne99 : in hex_char;
			correspondence_X51 : in hex_char;
			D05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_6;
	component railwaySignal_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R79_command : in routeCommands;
			R66_command : in routeCommands;
			--Ocupation level 0
			track_ne65 : in hex_char;
			correspondence_C119 : out hex_char;
			--Ocupation level 1
			track_ne992 : in hex_char;
			correspondence_J40 : in hex_char;
			Sw01_state : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			correspondence_L31 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_7;
	component railwaySignal_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R57_command : in routeCommands;
			R58_command : in routeCommands;
			R38_command : in routeCommands;
			--Ocupation level 0
			track_ne910 : in hex_char;
			correspondence_S81 : out hex_char;
			--Ocupation level 1
			track_ne130 : in hex_char;
			track_ne135 : in hex_char;
			correspondence_S107 : in hex_char;
			correspondence_B80 : in hex_char;
			D10_state : in hex_char;
			--Ocupation level 2
			track_ne129 : in hex_char;
			track_ne450 : in hex_char;
			track_ne114 : in hex_char;
			track_ne127 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_T07 : in hex_char;
			correspondence_S104 : in hex_char;
			D23_state : in hex_char;
			D12_state : in hex_char;
			D24_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_8;
	component railwaySignal_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R26_command : in routeCommands;
			R8_command : in routeCommands;
			R28_command : in routeCommands;
			--Ocupation level 0
			track_ne912 : in hex_char;
			correspondence_J45 : out hex_char;
			--Ocupation level 1
			track_ne101 : in hex_char;
			correspondence_J43 : in hex_char;
			D09_state : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			correspondence_X53 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_9;
	component railwaySignal_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			R37_command : in routeCommands;
			--Ocupation level 0
			track_ne912 : in hex_char;
			correspondence_S110 : out hex_char;
			--Ocupation level 1
			track_ne131 : in hex_char;
			track_ne465 : in hex_char;
			track_ne132 : in hex_char;
			correspondence_T09 : in hex_char;
			correspondence_J46 : in hex_char;
			D20_state : in hex_char;
			D21_state : in hex_char;
			--Ocupation level 2
			track_ne114 : in hex_char;
			correspondence_L29 : in hex_char;
			D23_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_10;
	component railwaySignal_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R17_command : in routeCommands;
			R27_command : in routeCommands;
			R71_command : in routeCommands;
			R73_command : in routeCommands;
			--Ocupation level 0
			track_ne114 : in hex_char;
			correspondence_L29 : out hex_char;
			correspondence_J48 : in hex_char;
			--Ocupation level 2
			track_ne102 : in hex_char;
			correspondence_T11 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_11;
	component railwaySignal_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R29_command : in routeCommands;
			R17_command : in routeCommands;
			--Ocupation level 0
			track_ne114 : in hex_char;
			correspondence_J48 : out hex_char;
			--Ocupation level 1
			track_ne102 : in hex_char;
			correspondence_T11 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_12;
	component railwaySignal_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R10_command : in routeCommands;
			--Ocupation level 0
			track_ne114 : in hex_char;
			correspondence_S101 : out hex_char;
			--Ocupation level 1
			track_ne132 : in hex_char;
			track_ne129 : in hex_char;
			track_ne127 : in hex_char;
			track_ne130 : in hex_char;
			correspondence_J47 : in hex_char;
			correspondence_S117 : in hex_char;
			correspondence_C79 : in hex_char;
			D23_state : in hex_char;
			D12_state : in hex_char;
			--Ocupation level 2
			track_ne912 : in hex_char;
			track_ne910 : in hex_char;
			track_ne134 : in hex_char;
			track_ne135 : in hex_char;
			track_ne101 : in hex_char;
			correspondence_J45 : in hex_char;
			correspondence_J43 : in hex_char;
			correspondence_T23 : in hex_char;
			D20_state : in hex_char;
			D09_state : in hex_char;
			D10_state : in hex_char;
			D24_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_13;
	component railwaySignal_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			R39_command : in routeCommands;
			--Ocupation level 0
			track_ne288 : in hex_char;
			correspondence_S69 : out hex_char;
			--Ocupation level 1
			track_ne295 : in hex_char;
			track_ne110 : in hex_char;
			correspondence_C70 : in hex_char;
			correspondence_B68 : in hex_char;
			D03_state : in hex_char;
			--Ocupation level 2
			track_ne297 : in hex_char;
			track_ne384 : in hex_char;
			correspondence_S126 : in hex_char;
			D04_state : in hex_char;
			Sw02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_14;
	component railwaySignal_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R20_command : in routeCommands;
			R2_command : in routeCommands;
			R22_command : in routeCommands;
			--Ocupation level 0
			track_ne290 : in hex_char;
			correspondence_J35 : out hex_char;
			--Ocupation level 1
			track_ne991 : in hex_char;
			correspondence_T01 : in hex_char;
			D01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_15;
	component railwaySignal_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			R40_command : in routeCommands;
			--Ocupation level 0
			track_ne290 : in hex_char;
			correspondence_S86 : out hex_char;
			--Ocupation level 1
			track_ne292 : in hex_char;
			track_ne111 : in hex_char;
			track_ne377 : in hex_char;
			correspondence_J36 : in hex_char;
			correspondence_T03 : in hex_char;
			D14_state : in hex_char;
			D15_state : in hex_char;
			--Ocupation level 2
			track_ne996 : in hex_char;
			correspondence_J38 : in hex_char;
			Sw04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_16;
	component railwaySignal_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R21_command : in routeCommands;
			R61_command : in routeCommands;
			--Ocupation level 0
			track_ne292 : in hex_char;
			correspondence_J36 : out hex_char;
			--Ocupation level 1
			track_ne996 : in hex_char;
			correspondence_J38 : in hex_char;
			Sw04_state : in hex_char;
			--Ocupation level 2
			track_ne98 : in hex_char;
			correspondence_L30 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_17;
	component railwaySignal_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R22_command : in routeCommands;
			R88_command : in routeCommands;
			--Ocupation level 0
			track_ne292 : in hex_char;
			correspondence_J37 : out hex_char;
			--Ocupation level 1
			track_ne290 : in hex_char;
			correspondence_J35 : in hex_char;
			D14_state : in hex_char;
			--Ocupation level 2
			track_ne991 : in hex_char;
			correspondence_T01 : in hex_char;
			D01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_18;
	component railwaySignal_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R41_command : in routeCommands;
			R46_command : in routeCommands;
			--Ocupation level 0
			track_ne295 : in hex_char;
			correspondence_C67 : out hex_char;
			--Ocupation level 1
			track_ne288 : in hex_char;
			track_ne991 : in hex_char;
			correspondence_T01 : in hex_char;
			D01_state : in hex_char;
			D03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_19;
	component railwaySignal_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R45_command : in routeCommands;
			R43_command : in routeCommands;
			--Ocupation level 0
			track_ne295 : in hex_char;
			correspondence_C70 : out hex_char;
			--Ocupation level 1
			track_ne297 : in hex_char;
			correspondence_S126 : in hex_char;
			D04_state : in hex_char;
			--Ocupation level 2
			track_ne996 : in hex_char;
			track_ne997 : in hex_char;
			track_ne995 : in hex_char;
			correspondence_T27 : in hex_char;
			correspondence_J38 : in hex_char;
			Sw03_state : in hex_char;
			Sw04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_20;
	component railwaySignal_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			R85_command : in routeCommands;
			R89_command : in routeCommands;
			--Ocupation level 0
			track_ne297 : in hex_char;
			correspondence_S71 : out hex_char;
			--Ocupation level 1
			track_ne295 : in hex_char;
			track_ne384 : in hex_char;
			correspondence_C67 : in hex_char;
			correspondence_S84 : in hex_char;
			D04_state : in hex_char;
			--Ocupation level 2
			track_ne991 : in hex_char;
			track_ne288 : in hex_char;
			track_ne104 : in hex_char;
			track_ne110 : in hex_char;
			correspondence_T01 : in hex_char;
			correspondence_T13 : in hex_char;
			D01_state : in hex_char;
			D03_state : in hex_char;
			Sw02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_21;
	component railwaySignal_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R86_command : in routeCommands;
			R87_command : in routeCommands;
			R11_command : in routeCommands;
			R42_command : in routeCommands;
			R45_command : in routeCommands;
			--Ocupation level 0
			track_ne297 : in hex_char;
			correspondence_S126 : out hex_char;
			--Ocupation level 1
			track_ne995 : in hex_char;
			track_ne997 : in hex_char;
			track_ne996 : in hex_char;
			correspondence_T27 : in hex_char;
			correspondence_J38 : in hex_char;
			Sw03_state : in hex_char;
			Sw04_state : in hex_char;
			--Ocupation level 2
			track_ne98 : in hex_char;
			correspondence_L30 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_22;
	component railwaySignal_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R12_command : in routeCommands;
			R62_command : in routeCommands;
			--Ocupation level 0
			track_ne377 : in hex_char;
			correspondence_T03 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_23;
	component railwaySignal_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R2_command : in routeCommands;
			R3_command : in routeCommands;
			--Ocupation level 0
			track_ne377 : in hex_char;
			correspondence_T04 : out hex_char;
			--Ocupation level 1
			track_ne111 : in hex_char;
			track_ne290 : in hex_char;
			track_ne113 : in hex_char;
			correspondence_J35 : in hex_char;
			correspondence_T15 : in hex_char;
			D14_state : in hex_char;
			D15_state : in hex_char;
			--Ocupation level 2
			track_ne991 : in hex_char;
			correspondence_T01 : in hex_char;
			D01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_24;
	component railwaySignal_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R59_command : in routeCommands;
			R60_command : in routeCommands;
			R47_command : in routeCommands;
			--Ocupation level 0
			track_ne384 : in hex_char;
			correspondence_S84 : out hex_char;
			--Ocupation level 1
			track_ne104 : in hex_char;
			track_ne110 : in hex_char;
			track_ne288 : in hex_char;
			track_ne991 : in hex_char;
			correspondence_T13 : in hex_char;
			correspondence_T01 : in hex_char;
			Sw02_state : in hex_char;
			D01_state : in hex_char;
			D03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_25;
	component railwaySignal_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			R81_command : in routeCommands;
			R82_command : in routeCommands;
			--Ocupation level 0
			track_ne400 : in hex_char;
			correspondence_S74 : out hex_char;
			--Ocupation level 1
			track_ne404 : in hex_char;
			track_ne407 : in hex_char;
			correspondence_C76 : in hex_char;
			correspondence_S93 : in hex_char;
			D07_state : in hex_char;
			--Ocupation level 2
			track_ne61 : in hex_char;
			track_ne98 : in hex_char;
			track_ne99 : in hex_char;
			track_ne122 : in hex_char;
			track_ne123 : in hex_char;
			correspondence_X51 : in hex_char;
			correspondence_T17 : in hex_char;
			D05_state : in hex_char;
			D08_state : in hex_char;
			D16_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_26;
	component railwaySignal_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R83_command : in routeCommands;
			R84_command : in routeCommands;
			R13_command : in routeCommands;
			R48_command : in routeCommands;
			R52_command : in routeCommands;
			--Ocupation level 0
			track_ne400 : in hex_char;
			correspondence_S123 : out hex_char;
			--Ocupation level 1
			track_ne993 : in hex_char;
			track_ne994 : in hex_char;
			track_ne992 : in hex_char;
			correspondence_T25 : in hex_char;
			correspondence_J40 : in hex_char;
			Sw05_state : in hex_char;
			Sw01_state : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			correspondence_L31 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_27;
	component railwaySignal_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R48_command : in routeCommands;
			R53_command : in routeCommands;
			--Ocupation level 0
			track_ne404 : in hex_char;
			correspondence_C73 : out hex_char;
			--Ocupation level 1
			track_ne400 : in hex_char;
			correspondence_S123 : in hex_char;
			D07_state : in hex_char;
			--Ocupation level 2
			track_ne994 : in hex_char;
			track_ne992 : in hex_char;
			track_ne993 : in hex_char;
			correspondence_T25 : in hex_char;
			correspondence_J40 : in hex_char;
			Sw05_state : in hex_char;
			Sw01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_28;
	component railwaySignal_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R51_command : in routeCommands;
			R49_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne404 : in hex_char;
			correspondence_C76 : out hex_char;
			--Ocupation level 1
			track_ne61 : in hex_char;
			track_ne99 : in hex_char;
			track_ne98 : in hex_char;
			correspondence_X51 : in hex_char;
			D05_state : in hex_char;
			D08_state : in hex_char;
			--Ocupation level 2
			track_ne996 : in hex_char;
			correspondence_S129 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_29;
	component railwaySignal_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			R50_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne407 : in hex_char;
			correspondence_S93 : out hex_char;
			--Ocupation level 1
			track_ne122 : in hex_char;
			track_ne123 : in hex_char;
			track_ne61 : in hex_char;
			track_ne99 : in hex_char;
			track_ne98 : in hex_char;
			correspondence_T17 : in hex_char;
			correspondence_X51 : in hex_char;
			D16_state : in hex_char;
			D05_state : in hex_char;
			D08_state : in hex_char;
			--Ocupation level 2
			track_ne996 : in hex_char;
			correspondence_S129 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_30;
	component railwaySignal_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R14_command : in routeCommands;
			R67_command : in routeCommands;
			--Ocupation level 0
			track_ne421 : in hex_char;
			correspondence_T05 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_31;
	component railwaySignal_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			R5_command : in routeCommands;
			--Ocupation level 0
			track_ne421 : in hex_char;
			correspondence_T06 : out hex_char;
			--Ocupation level 1
			track_ne124 : in hex_char;
			track_ne63 : in hex_char;
			track_ne126 : in hex_char;
			correspondence_C54 : in hex_char;
			correspondence_T19 : in hex_char;
			D18_state : in hex_char;
			D19_state : in hex_char;
			--Ocupation level 2
			track_ne98 : in hex_char;
			track_ne99 : in hex_char;
			correspondence_X51 : in hex_char;
			D05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_32;
	component railwaySignal_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R72_command : in routeCommands;
			R74_command : in routeCommands;
			--Ocupation level 0
			track_ne450 : in hex_char;
			correspondence_T07 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_33;
	component railwaySignal_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R6_command : in routeCommands;
			R7_command : in routeCommands;
			--Ocupation level 0
			track_ne450 : in hex_char;
			correspondence_T08 : out hex_char;
			--Ocupation level 1
			track_ne127 : in hex_char;
			track_ne130 : in hex_char;
			correspondence_S117 : in hex_char;
			correspondence_C79 : in hex_char;
			D12_state : in hex_char;
			--Ocupation level 2
			track_ne910 : in hex_char;
			track_ne134 : in hex_char;
			track_ne135 : in hex_char;
			track_ne101 : in hex_char;
			correspondence_J43 : in hex_char;
			correspondence_T23 : in hex_char;
			D09_state : in hex_char;
			D10_state : in hex_char;
			D24_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_34;
	component railwaySignal_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R15_command : in routeCommands;
			R75_command : in routeCommands;
			--Ocupation level 0
			track_ne465 : in hex_char;
			correspondence_T09 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_35;
	component railwaySignal_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R8_command : in routeCommands;
			R9_command : in routeCommands;
			--Ocupation level 0
			track_ne465 : in hex_char;
			correspondence_T10 : out hex_char;
			--Ocupation level 1
			track_ne131 : in hex_char;
			track_ne912 : in hex_char;
			track_ne133 : in hex_char;
			correspondence_J45 : in hex_char;
			correspondence_T21 : in hex_char;
			D20_state : in hex_char;
			D21_state : in hex_char;
			--Ocupation level 2
			track_ne101 : in hex_char;
			correspondence_J43 : in hex_char;
			D09_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_36;
	component railwaySignal_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R18_command : in routeCommands;
			R23_command : in routeCommands;
			--Ocupation level 0
			track_ne98 : in hex_char;
			correspondence_L30 : out hex_char;
			correspondence_X50 : in hex_char;
			--Ocupation level 2
			track_ne99 : in hex_char;
			correspondence_S55 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_37;
	component railwaySignal_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R30_command : in routeCommands;
			R18_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne98 : in hex_char;
			correspondence_X50 : out hex_char;
			--Ocupation level 1
			track_ne99 : in hex_char;
			correspondence_S55 : in hex_char;
			--Ocupation level 2
			track_ne63 : in hex_char;
			track_ne61 : in hex_char;
			correspondence_S78 : in hex_char;
			correspondence_S95 : in hex_char;
			D05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_38;
	component railwaySignal_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R31_command : in routeCommands;
			R34_command : in routeCommands;
			R51_command : in routeCommands;
			R64_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne98 : in hex_char;
			correspondence_X51 : out hex_char;
			--Ocupation level 1
			track_ne996 : in hex_char;
			correspondence_S129 : in hex_char;
			--Ocupation level 2
			track_ne292 : in hex_char;
			track_ne997 : in hex_char;
			track_ne297 : in hex_char;
			correspondence_J37 : in hex_char;
			correspondence_S71 : in hex_char;
			Sw04_state : in hex_char;
			Sw03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_39;
	component railwaySignal_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R35_command : in routeCommands;
			R36_command : in routeCommands;
			R30_command : in routeCommands;
			--Ocupation level 0
			track_ne99 : in hex_char;
			correspondence_S55 : out hex_char;
			--Ocupation level 1
			track_ne61 : in hex_char;
			track_ne63 : in hex_char;
			correspondence_S78 : in hex_char;
			correspondence_S95 : in hex_char;
			D05_state : in hex_char;
			--Ocupation level 2
			track_ne404 : in hex_char;
			track_ne123 : in hex_char;
			track_ne421 : in hex_char;
			track_ne65 : in hex_char;
			track_ne124 : in hex_char;
			correspondence_C73 : in hex_char;
			correspondence_B77 : in hex_char;
			correspondence_C119 : in hex_char;
			correspondence_T05 : in hex_char;
			D08_state : in hex_char;
			D18_state : in hex_char;
			D19_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_40;
	component railwaySignal_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R19_command : in routeCommands;
			R24_command : in routeCommands;
			--Ocupation level 0
			track_ne100 : in hex_char;
			correspondence_L31 : out hex_char;
			correspondence_X52 : in hex_char;
			--Ocupation level 2
			track_ne101 : in hex_char;
			correspondence_S59 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_41;
	component railwaySignal_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R32_command : in routeCommands;
			R19_command : in routeCommands;
			Lc04_state : in hex_char;
			--Ocupation level 0
			track_ne100 : in hex_char;
			correspondence_X52 : out hex_char;
			--Ocupation level 1
			track_ne101 : in hex_char;
			correspondence_S59 : in hex_char;
			--Ocupation level 2
			track_ne910 : in hex_char;
			track_ne912 : in hex_char;
			correspondence_S110 : in hex_char;
			correspondence_S81 : in hex_char;
			D09_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_42;
	component railwaySignal_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R33_command : in routeCommands;
			R25_command : in routeCommands;
			Lc04_state : in hex_char;
			--Ocupation level 0
			track_ne100 : in hex_char;
			correspondence_X53 : out hex_char;
			--Ocupation level 1
			track_ne992 : in hex_char;
			correspondence_S120 : in hex_char;
			--Ocupation level 2
			track_ne994 : in hex_char;
			track_ne65 : in hex_char;
			track_ne400 : in hex_char;
			correspondence_C94 : in hex_char;
			correspondence_S74 : in hex_char;
			Sw01_state : in hex_char;
			Sw05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_43;
	component railwaySignal_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			R55_command : in routeCommands;
			R77_command : in routeCommands;
			--Ocupation level 0
			track_ne101 : in hex_char;
			correspondence_J43 : out hex_char;
			--Ocupation level 1
			track_ne100 : in hex_char;
			correspondence_X53 : in hex_char;
			--Ocupation level 2
			track_ne992 : in hex_char;
			correspondence_S120 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_44;
	component railwaySignal_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R37_command : in routeCommands;
			R38_command : in routeCommands;
			R32_command : in routeCommands;
			--Ocupation level 0
			track_ne101 : in hex_char;
			correspondence_S59 : out hex_char;
			--Ocupation level 1
			track_ne912 : in hex_char;
			track_ne910 : in hex_char;
			correspondence_S110 : in hex_char;
			correspondence_S81 : in hex_char;
			D09_state : in hex_char;
			--Ocupation level 2
			track_ne131 : in hex_char;
			track_ne132 : in hex_char;
			track_ne465 : in hex_char;
			track_ne130 : in hex_char;
			track_ne135 : in hex_char;
			correspondence_T09 : in hex_char;
			correspondence_J46 : in hex_char;
			correspondence_S107 : in hex_char;
			correspondence_B80 : in hex_char;
			D20_state : in hex_char;
			D21_state : in hex_char;
			D10_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_45;
	component railwaySignal_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R29_command : in routeCommands;
			--Ocupation level 0
			track_ne102 : in hex_char;
			correspondence_T11 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_46;
	component railwaySignal_47 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R10_command : in routeCommands;
			--Ocupation level 0
			track_ne102 : in hex_char;
			correspondence_T12 : out hex_char;
			--Ocupation level 1
			track_ne114 : in hex_char;
			correspondence_S101 : in hex_char;
			--Ocupation level 2
			track_ne130 : in hex_char;
			track_ne129 : in hex_char;
			track_ne132 : in hex_char;
			track_ne127 : in hex_char;
			correspondence_J47 : in hex_char;
			correspondence_S117 : in hex_char;
			correspondence_C79 : in hex_char;
			D23_state : in hex_char;
			D12_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_47;
	component railwaySignal_48 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R59_command : in routeCommands;
			--Ocupation level 0
			track_ne104 : in hex_char;
			correspondence_T13 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_48;
	component railwaySignal_49 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R11_command : in routeCommands;
			--Ocupation level 0
			track_ne104 : in hex_char;
			correspondence_T14 : out hex_char;
			--Ocupation level 1
			track_ne384 : in hex_char;
			track_ne297 : in hex_char;
			correspondence_S126 : in hex_char;
			D04_state : in hex_char;
			Sw02_state : in hex_char;
			--Ocupation level 2
			track_ne996 : in hex_char;
			track_ne997 : in hex_char;
			track_ne995 : in hex_char;
			correspondence_T27 : in hex_char;
			correspondence_J38 : in hex_char;
			Sw03_state : in hex_char;
			Sw04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_49;
	component railwaySignal_50 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			--Ocupation level 0
			track_ne110 : in hex_char;
			correspondence_B68 : out hex_char;
			--Ocupation level 1
			track_ne384 : in hex_char;
			track_ne297 : in hex_char;
			correspondence_S126 : in hex_char;
			D04_state : in hex_char;
			Sw02_state : in hex_char;
			--Ocupation level 2
			track_ne996 : in hex_char;
			track_ne997 : in hex_char;
			track_ne995 : in hex_char;
			correspondence_T27 : in hex_char;
			correspondence_J38 : in hex_char;
			Sw03_state : in hex_char;
			Sw04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_50;
	component railwaySignal_51 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R3_command : in routeCommands;
			--Ocupation level 0
			track_ne113 : in hex_char;
			correspondence_T15 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_51;
	component railwaySignal_52 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R12_command : in routeCommands;
			--Ocupation level 0
			track_ne113 : in hex_char;
			correspondence_T16 : out hex_char;
			--Ocupation level 1
			track_ne377 : in hex_char;
			correspondence_T03 : in hex_char;
			D15_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_52;
	component railwaySignal_53 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R63_command : in routeCommands;
			--Ocupation level 0
			track_ne122 : in hex_char;
			correspondence_T17 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_53;
	component railwaySignal_54 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R13_command : in routeCommands;
			--Ocupation level 0
			track_ne122 : in hex_char;
			correspondence_T18 : out hex_char;
			--Ocupation level 1
			track_ne407 : in hex_char;
			track_ne400 : in hex_char;
			correspondence_S123 : in hex_char;
			D07_state : in hex_char;
			D16_state : in hex_char;
			--Ocupation level 2
			track_ne994 : in hex_char;
			track_ne992 : in hex_char;
			track_ne993 : in hex_char;
			correspondence_T25 : in hex_char;
			correspondence_J40 : in hex_char;
			Sw05_state : in hex_char;
			Sw01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_54;
	component railwaySignal_55 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R52_command : in routeCommands;
			R54_command : in routeCommands;
			--Ocupation level 0
			track_ne123 : in hex_char;
			correspondence_B77 : out hex_char;
			--Ocupation level 1
			track_ne407 : in hex_char;
			track_ne400 : in hex_char;
			correspondence_S123 : in hex_char;
			D07_state : in hex_char;
			D16_state : in hex_char;
			--Ocupation level 2
			track_ne994 : in hex_char;
			track_ne992 : in hex_char;
			track_ne993 : in hex_char;
			correspondence_T25 : in hex_char;
			correspondence_J40 : in hex_char;
			Sw05_state : in hex_char;
			Sw01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_55;
	component railwaySignal_56 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R5_command : in routeCommands;
			--Ocupation level 0
			track_ne126 : in hex_char;
			correspondence_T19 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_56;
	component railwaySignal_57 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R14_command : in routeCommands;
			--Ocupation level 0
			track_ne126 : in hex_char;
			correspondence_T20 : out hex_char;
			--Ocupation level 1
			track_ne421 : in hex_char;
			correspondence_T05 : in hex_char;
			D19_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_57;
	component railwaySignal_58 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			R16_command : in routeCommands;
			R56_command : in routeCommands;
			--Ocupation level 0
			track_ne127 : in hex_char;
			correspondence_S104 : out hex_char;
			--Ocupation level 1
			track_ne129 : in hex_char;
			track_ne114 : in hex_char;
			track_ne450 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_T07 : in hex_char;
			D23_state : in hex_char;
			D12_state : in hex_char;
			correspondence_J48 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_58;
	component railwaySignal_59 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			R6_command : in routeCommands;
			R69_command : in routeCommands;
			--Ocupation level 0
			track_ne127 : in hex_char;
			correspondence_S117 : out hex_char;
			--Ocupation level 1
			track_ne135 : in hex_char;
			track_ne910 : in hex_char;
			track_ne101 : in hex_char;
			track_ne134 : in hex_char;
			correspondence_J43 : in hex_char;
			correspondence_T23 : in hex_char;
			D09_state : in hex_char;
			D10_state : in hex_char;
			D24_state : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			correspondence_X53 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_59;
	component railwaySignal_60 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R55_command : in routeCommands;
			R7_command : in routeCommands;
			R70_command : in routeCommands;
			--Ocupation level 0
			track_ne130 : in hex_char;
			correspondence_C79 : out hex_char;
			--Ocupation level 1
			track_ne910 : in hex_char;
			track_ne101 : in hex_char;
			correspondence_J43 : in hex_char;
			D09_state : in hex_char;
			D10_state : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			correspondence_X53 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_60;
	component railwaySignal_61 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			R57_command : in routeCommands;
			--Ocupation level 0
			track_ne130 : in hex_char;
			correspondence_S107 : out hex_char;
			--Ocupation level 1
			track_ne129 : in hex_char;
			track_ne114 : in hex_char;
			track_ne450 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_T07 : in hex_char;
			D23_state : in hex_char;
			D12_state : in hex_char;
			correspondence_J48 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_61;
	component railwaySignal_62 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R27_command : in routeCommands;
			R76_command : in routeCommands;
			--Ocupation level 0
			track_ne132 : in hex_char;
			correspondence_J46 : out hex_char;
			--Ocupation level 1
			track_ne114 : in hex_char;
			correspondence_L29 : in hex_char;
			D23_state : in hex_char;
			correspondence_J48 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_62;
	component railwaySignal_63 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R28_command : in routeCommands;
			R68_command : in routeCommands;
			--Ocupation level 0
			track_ne132 : in hex_char;
			correspondence_J47 : out hex_char;
			--Ocupation level 1
			track_ne912 : in hex_char;
			correspondence_J45 : in hex_char;
			D20_state : in hex_char;
			--Ocupation level 2
			track_ne101 : in hex_char;
			correspondence_J43 : in hex_char;
			D09_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_63;
	component railwaySignal_64 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R9_command : in routeCommands;
			--Ocupation level 0
			track_ne133 : in hex_char;
			correspondence_T21 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_64;
	component railwaySignal_65 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R15_command : in routeCommands;
			--Ocupation level 0
			track_ne133 : in hex_char;
			correspondence_T22 : out hex_char;
			--Ocupation level 1
			track_ne465 : in hex_char;
			correspondence_T09 : in hex_char;
			D21_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_65;
	component railwaySignal_66 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R78_command : in routeCommands;
			--Ocupation level 0
			track_ne134 : in hex_char;
			correspondence_T23 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_66;
	component railwaySignal_67 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R16_command : in routeCommands;
			--Ocupation level 0
			track_ne134 : in hex_char;
			correspondence_T24 : out hex_char;
			--Ocupation level 1
			track_ne127 : in hex_char;
			correspondence_S104 : in hex_char;
			D24_state : in hex_char;
			--Ocupation level 2
			track_ne129 : in hex_char;
			track_ne450 : in hex_char;
			track_ne114 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_T07 : in hex_char;
			D23_state : in hex_char;
			D12_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_67;
	component railwaySignal_68 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			--Ocupation level 0
			track_ne135 : in hex_char;
			correspondence_B80 : out hex_char;
			--Ocupation level 1
			track_ne127 : in hex_char;
			correspondence_S104 : in hex_char;
			D24_state : in hex_char;
			--Ocupation level 2
			track_ne129 : in hex_char;
			track_ne450 : in hex_char;
			track_ne114 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_T07 : in hex_char;
			D23_state : in hex_char;
			D12_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_68;
	component railwaySignal_69 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R24_command : in routeCommands;
			R79_command : in routeCommands;
			R84_command : in routeCommands;
			--Ocupation level 0
			track_ne992 : in hex_char;
			correspondence_J40 : out hex_char;
			--Ocupation level 1
			track_ne100 : in hex_char;
			correspondence_L31 : in hex_char;
			correspondence_X52 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_69;
	component railwaySignal_70 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R80_command : in routeCommands;
			R81_command : in routeCommands;
			R33_command : in routeCommands;
			--Ocupation level 0
			track_ne992 : in hex_char;
			correspondence_S120 : out hex_char;
			--Ocupation level 1
			track_ne65 : in hex_char;
			track_ne994 : in hex_char;
			track_ne400 : in hex_char;
			correspondence_C94 : in hex_char;
			correspondence_S74 : in hex_char;
			Sw01_state : in hex_char;
			Sw05_state : in hex_char;
			--Ocupation level 2
			track_ne63 : in hex_char;
			track_ne407 : in hex_char;
			track_ne404 : in hex_char;
			correspondence_C54 : in hex_char;
			correspondence_C76 : in hex_char;
			correspondence_S93 : in hex_char;
			D18_state : in hex_char;
			D07_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_70;
	component railwaySignal_71 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R83_command : in routeCommands;
			--Ocupation level 0
			track_ne993 : in hex_char;
			correspondence_T25 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_71;
	component railwaySignal_72 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R82_command : in routeCommands;
			--Ocupation level 0
			track_ne993 : in hex_char;
			correspondence_C122 : out hex_char;
			--Ocupation level 1
			track_ne400 : in hex_char;
			correspondence_S74 : in hex_char;
			Sw05_state : in hex_char;
			--Ocupation level 2
			track_ne407 : in hex_char;
			track_ne404 : in hex_char;
			correspondence_C76 : in hex_char;
			correspondence_S93 : in hex_char;
			D07_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_72;
	component railwaySignal_73 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R86_command : in routeCommands;
			--Ocupation level 0
			track_ne995 : in hex_char;
			correspondence_T27 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_73;
	component railwaySignal_74 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R85_command : in routeCommands;
			--Ocupation level 0
			track_ne995 : in hex_char;
			correspondence_C125 : out hex_char;
			--Ocupation level 1
			track_ne297 : in hex_char;
			correspondence_S71 : in hex_char;
			Sw03_state : in hex_char;
			--Ocupation level 2
			track_ne384 : in hex_char;
			track_ne295 : in hex_char;
			correspondence_C67 : in hex_char;
			correspondence_S84 : in hex_char;
			D04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_74;
	component railwaySignal_75 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R23_command : in routeCommands;
			R21_command : in routeCommands;
			R87_command : in routeCommands;
			--Ocupation level 0
			track_ne996 : in hex_char;
			correspondence_J38 : out hex_char;
			--Ocupation level 1
			track_ne98 : in hex_char;
			correspondence_L30 : in hex_char;
			correspondence_X50 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_75;
	component railwaySignal_76 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R88_command : in routeCommands;
			R89_command : in routeCommands;
			R31_command : in routeCommands;
			--Ocupation level 0
			track_ne996 : in hex_char;
			correspondence_S129 : out hex_char;
			--Ocupation level 1
			track_ne292 : in hex_char;
			track_ne997 : in hex_char;
			track_ne297 : in hex_char;
			correspondence_J37 : in hex_char;
			correspondence_S71 : in hex_char;
			Sw04_state : in hex_char;
			Sw03_state : in hex_char;
			--Ocupation level 2
			track_ne290 : in hex_char;
			track_ne384 : in hex_char;
			track_ne295 : in hex_char;
			correspondence_J35 : in hex_char;
			correspondence_C67 : in hex_char;
			correspondence_S84 : in hex_char;
			D14_state : in hex_char;
			D04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_76;
	component node_0 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R1_command : in routeCommands;
			R20_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			R41_command : in routeCommands;
			R60_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_0;
	component node_1 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R35_command : in routeCommands;
			R51_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R64_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_1;
	component node_2 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R4_command : in routeCommands;
			R34_command : in routeCommands;
			R36_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R67_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_2;
	component node_3 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_3;
	component node_4 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R38_command : in routeCommands;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			R58_command : in routeCommands;
			R77_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_4;
	component node_5 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R8_command : in routeCommands;
			R26_command : in routeCommands;
			R28_command : in routeCommands;
			R37_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_5;
	component node_6 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R10_command : in routeCommands;
			R17_command : in routeCommands;
			R27_command : in routeCommands;
			R29_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R73_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_6;
	component node_7 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R39_command : in routeCommands;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			R60_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_7;
	component node_8 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R2_command : in routeCommands;
			R20_command : in routeCommands;
			R22_command : in routeCommands;
			R40_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_8;
	component node_9 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R21_command : in routeCommands;
			R22_command : in routeCommands;
			R61_command : in routeCommands;
			R88_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_9;
	component node_10 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R45_command : in routeCommands;
			R46_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_10;
	component node_11 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R11_command : in routeCommands;
			R42_command : in routeCommands;
			R45_command : in routeCommands;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			R87_command : in routeCommands;
			R89_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_11;
	component node_12 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R2_command : in routeCommands;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			R62_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_12;
	component node_13 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R11_command : in routeCommands;
			R42_command : in routeCommands;
			R47_command : in routeCommands;
			R59_command : in routeCommands;
			R60_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_13;
	component node_14 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R13_command : in routeCommands;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			R52_command : in routeCommands;
			R81_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			R84_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_14;
	component node_15 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R51_command : in routeCommands;
			R53_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_15;
	component node_16 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R13_command : in routeCommands;
			R50_command : in routeCommands;
			R52_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_16;
	component node_17 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R4_command : in routeCommands;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			R67_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_17;
	component node_18 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R6_command : in routeCommands;
			R7_command : in routeCommands;
			R72_command : in routeCommands;
			R74_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_18;
	component node_19 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R8_command : in routeCommands;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			R75_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_19;
	component node_20 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R18_command : in routeCommands;
			R23_command : in routeCommands;
			R30_command : in routeCommands;
			R31_command : in routeCommands;
			R34_command : in routeCommands;
			R51_command : in routeCommands;
			R64_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_20;
	component node_21 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R30_command : in routeCommands;
			R34_command : in routeCommands;
			R35_command : in routeCommands;
			R36_command : in routeCommands;
			R51_command : in routeCommands;
			R64_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_21;
	component node_22 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R19_command : in routeCommands;
			R24_command : in routeCommands;
			R25_command : in routeCommands;
			R32_command : in routeCommands;
			R33_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_22;
	component node_23 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			R32_command : in routeCommands;
			R37_command : in routeCommands;
			R38_command : in routeCommands;
			R55_command : in routeCommands;
			R77_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_23;
	component node_24 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R10_command : in routeCommands;
			R29_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_24;
	component node_25 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R11_command : in routeCommands;
			R59_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_25;
	component node_26 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			R60_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_26;
	component node_27 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R2_command : in routeCommands;
			R62_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_27;
	component node_28 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_28;
	component node_29 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R13_command : in routeCommands;
			R63_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_29;
	component node_30 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R52_command : in routeCommands;
			R54_command : in routeCommands;
			R64_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_30;
	component node_31 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R4_command : in routeCommands;
			R67_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_31;
	component node_32 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_32;
	component node_33 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R6_command : in routeCommands;
			R16_command : in routeCommands;
			R56_command : in routeCommands;
			R69_command : in routeCommands;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_33;
	component node_34 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R73_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_34;
	component node_35 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R7_command : in routeCommands;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			R70_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_35;
	component node_36 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R8_command : in routeCommands;
			R75_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_36;
	component node_37 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R27_command : in routeCommands;
			R28_command : in routeCommands;
			R68_command : in routeCommands;
			R76_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_37;
	component node_38 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_38;
	component node_39 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R16_command : in routeCommands;
			R78_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_39;
	component node_40 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R77_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_40;
	component node_41 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R24_command : in routeCommands;
			R33_command : in routeCommands;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			R81_command : in routeCommands;
			R84_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_41;
	component node_42 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_42;
	component node_43 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R81_command : in routeCommands;
			R84_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_43;
	component node_44 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_44;
	component node_45 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R21_command : in routeCommands;
			R23_command : in routeCommands;
			R31_command : in routeCommands;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			R89_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_45;
	component node_46 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R87_command : in routeCommands;
			R89_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_46;
--sw  R1 ['D01'] 
--dw  R1 [] 
--sc  R1 [] 
--lc  R1 [] 
	component route_0 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne991 : in hex_char;
			ne991_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			T02_state : in hex_char;
			T02_command : out routeCommands := RELEASE;
			S64_state : in hex_char;
			S64_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_0;
--sw  R2 ['D01', 'D14', 'D15'] 
--dw  R2 [] 
--sc  R2 [] 
--lc  R2 [] 
	component route_1 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne377 : in hex_char;
			ne377_command : out routeCommands := RELEASE;
			track_ne111 : in hex_char;
			ne111_command : out routeCommands := RELEASE;
			track_ne290 : in hex_char;
			ne290_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			D14_state : in hex_char;
			D14_command : out routeCommands := RELEASE;
			D15_state : in hex_char;
			D15_command : out routeCommands := RELEASE;
			T04_state : in hex_char;
			T04_command : out routeCommands := RELEASE;
			J35_state : in hex_char;
			J35_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_1;
--sw  R3 ['D15'] 
--dw  R3 [] 
--sc  R3 [] 
--lc  R3 [] 
	component route_2 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne377 : in hex_char;
			ne377_command : out routeCommands := RELEASE;
			track_ne113 : in hex_char;
			ne113_command : out routeCommands := RELEASE;
			D15_state : in hex_char;
			D15_command : out routeCommands := RELEASE;
			T04_state : in hex_char;
			T04_command : out routeCommands := RELEASE;
			T15_state : in hex_char;
			T15_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_2;
--sw  R4 ['D05', 'D18', 'D19'] 
--dw  R4 [] 
--sc  R4 [] 
--lc  R4 [] 
	component route_3 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne421 : in hex_char;
			ne421_command : out routeCommands := RELEASE;
			track_ne124 : in hex_char;
			ne124_command : out routeCommands := RELEASE;
			track_ne63 : in hex_char;
			ne63_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			D18_state : in hex_char;
			D18_command : out routeCommands := RELEASE;
			D19_state : in hex_char;
			D19_command : out routeCommands := RELEASE;
			T06_state : in hex_char;
			T06_command : out routeCommands := RELEASE;
			C54_state : in hex_char;
			C54_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_3;
--sw  R5 ['D19'] 
--dw  R5 [] 
--sc  R5 [] 
--lc  R5 [] 
	component route_4 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne421 : in hex_char;
			ne421_command : out routeCommands := RELEASE;
			track_ne126 : in hex_char;
			ne126_command : out routeCommands := RELEASE;
			D19_state : in hex_char;
			D19_command : out routeCommands := RELEASE;
			T06_state : in hex_char;
			T06_command : out routeCommands := RELEASE;
			T19_state : in hex_char;
			T19_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_4;
--sw  R6 ['D10', 'D09', 'D24'] 
--dw  R6 ['D12'] 
--sc  R6 [] 
--lc  R6 [] 
	component route_5 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne450 : in hex_char;
			ne450_command : out routeCommands := RELEASE;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D24_state : in hex_char;
			D24_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			T08_state : in hex_char;
			T08_command : out routeCommands := RELEASE;
			S117_state : in hex_char;
			S117_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_5;
--sw  R7 ['D10', 'D09'] 
--dw  R7 ['D12'] 
--sc  R7 [] 
--lc  R7 [] 
	component route_6 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne450 : in hex_char;
			ne450_command : out routeCommands := RELEASE;
			track_ne130 : in hex_char;
			ne130_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			T08_state : in hex_char;
			T08_command : out routeCommands := RELEASE;
			C79_state : in hex_char;
			C79_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_6;
--sw  R8 ['D09', 'D20', 'D21'] 
--dw  R8 [] 
--sc  R8 [] 
--lc  R8 [] 
	component route_7 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne465 : in hex_char;
			ne465_command : out routeCommands := RELEASE;
			track_ne131 : in hex_char;
			ne131_command : out routeCommands := RELEASE;
			track_ne912 : in hex_char;
			ne912_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D20_state : in hex_char;
			D20_command : out routeCommands := RELEASE;
			D21_state : in hex_char;
			D21_command : out routeCommands := RELEASE;
			T10_state : in hex_char;
			T10_command : out routeCommands := RELEASE;
			J45_state : in hex_char;
			J45_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_7;
--sw  R9 ['D21'] 
--dw  R9 [] 
--sc  R9 [] 
--lc  R9 [] 
	component route_8 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne465 : in hex_char;
			ne465_command : out routeCommands := RELEASE;
			track_ne133 : in hex_char;
			ne133_command : out routeCommands := RELEASE;
			D21_state : in hex_char;
			D21_command : out routeCommands := RELEASE;
			T10_state : in hex_char;
			T10_command : out routeCommands := RELEASE;
			T21_state : in hex_char;
			T21_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_8;
--sw  R10 ['D23'] 
--dw  R10 [] 
--sc  R10 [] 
--lc  R10 [] 
	component route_9 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne102 : in hex_char;
			ne102_command : out routeCommands := RELEASE;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			T12_state : in hex_char;
			T12_command : out routeCommands := RELEASE;
			S101_state : in hex_char;
			S101_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_9;
--sw  R11 ['D04', 'Sw03', 'Sw02'] 
--dw  R11 [] 
--sc  R11 [] 
--lc  R11 [] 
	component route_10 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne104 : in hex_char;
			ne104_command : out routeCommands := RELEASE;
			track_ne384 : in hex_char;
			ne384_command : out routeCommands := RELEASE;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			Sw02_state : in hex_char;
			Sw02_command : out routeCommands := RELEASE;
			T14_state : in hex_char;
			T14_command : out routeCommands := RELEASE;
			S126_state : in hex_char;
			S126_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_10;
--sw  R12 ['D15'] 
--dw  R12 [] 
--sc  R12 [] 
--lc  R12 [] 
	component route_11 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne113 : in hex_char;
			ne113_command : out routeCommands := RELEASE;
			track_ne377 : in hex_char;
			ne377_command : out routeCommands := RELEASE;
			D15_state : in hex_char;
			D15_command : out routeCommands := RELEASE;
			T16_state : in hex_char;
			T16_command : out routeCommands := RELEASE;
			T03_state : in hex_char;
			T03_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_11;
--sw  R13 ['D07', 'Sw05', 'D16'] 
--dw  R13 [] 
--sc  R13 [] 
--lc  R13 [] 
	component route_12 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne122 : in hex_char;
			ne122_command : out routeCommands := RELEASE;
			track_ne407 : in hex_char;
			ne407_command : out routeCommands := RELEASE;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			D16_state : in hex_char;
			D16_command : out routeCommands := RELEASE;
			T18_state : in hex_char;
			T18_command : out routeCommands := RELEASE;
			S123_state : in hex_char;
			S123_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_12;
--sw  R14 ['D19'] 
--dw  R14 [] 
--sc  R14 [] 
--lc  R14 [] 
	component route_13 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne126 : in hex_char;
			ne126_command : out routeCommands := RELEASE;
			track_ne421 : in hex_char;
			ne421_command : out routeCommands := RELEASE;
			D19_state : in hex_char;
			D19_command : out routeCommands := RELEASE;
			T20_state : in hex_char;
			T20_command : out routeCommands := RELEASE;
			T05_state : in hex_char;
			T05_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_13;
--sw  R15 ['D21'] 
--dw  R15 [] 
--sc  R15 [] 
--lc  R15 [] 
	component route_14 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne133 : in hex_char;
			ne133_command : out routeCommands := RELEASE;
			track_ne465 : in hex_char;
			ne465_command : out routeCommands := RELEASE;
			D21_state : in hex_char;
			D21_command : out routeCommands := RELEASE;
			T22_state : in hex_char;
			T22_command : out routeCommands := RELEASE;
			T09_state : in hex_char;
			T09_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_14;
--sw  R16 ['D23', 'D24'] 
--dw  R16 [] 
--sc  R16 [] 
--lc  R16 [] 
	component route_15 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne134 : in hex_char;
			ne134_command : out routeCommands := RELEASE;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			D24_state : in hex_char;
			D24_command : out routeCommands := RELEASE;
			T24_state : in hex_char;
			T24_command : out routeCommands := RELEASE;
			S104_state : in hex_char;
			S104_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_15;
--sw  R17 [] 
--dw  R17 [] 
--sc  R17 [] 
--lc  R17 [] 
	component route_16 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			L29_state : in hex_char;
			L29_command : out routeCommands := RELEASE;
			J48_state : in hex_char;
			J48_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_16;
--sw  R18 [] 
--dw  R18 [] 
--sc  R18 [] 
--lc  R18 [] 
	component route_17 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			L30_state : in hex_char;
			L30_command : out routeCommands := RELEASE;
			X50_state : in hex_char;
			X50_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_17;
--sw  R19 [] 
--dw  R19 [] 
--sc  R19 [] 
--lc  R19 [] 
	component route_18 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			L31_state : in hex_char;
			L31_command : out routeCommands := RELEASE;
			X52_state : in hex_char;
			X52_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_18;
--sw  R20 ['D01'] 
--dw  R20 [] 
--sc  R20 [] 
--lc  R20 [] 
	component route_19 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne290 : in hex_char;
			ne290_command : out routeCommands := RELEASE;
			track_ne991 : in hex_char;
			ne991_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			J35_state : in hex_char;
			J35_command : out routeCommands := RELEASE;
			T01_state : in hex_char;
			T01_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_19;
--sw  R21 ['Sw04'] 
--dw  R21 [] 
--sc  R21 [] 
--lc  R21 [] 
	component route_20 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne292 : in hex_char;
			ne292_command : out routeCommands := RELEASE;
			track_ne996 : in hex_char;
			ne996_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			J36_state : in hex_char;
			J36_command : out routeCommands := RELEASE;
			J38_state : in hex_char;
			J38_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_20;
--sw  R22 ['D01', 'D14'] 
--dw  R22 [] 
--sc  R22 [] 
--lc  R22 [] 
	component route_21 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne292 : in hex_char;
			ne292_command : out routeCommands := RELEASE;
			track_ne290 : in hex_char;
			ne290_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			D14_state : in hex_char;
			D14_command : out routeCommands := RELEASE;
			J37_state : in hex_char;
			J37_command : out routeCommands := RELEASE;
			J35_state : in hex_char;
			J35_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_21;
--sw  R23 [] 
--dw  R23 [] 
--sc  R23 [] 
--lc  R23 [] 
	component route_22 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne996 : in hex_char;
			ne996_command : out routeCommands := RELEASE;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			J38_state : in hex_char;
			J38_command : out routeCommands := RELEASE;
			L30_state : in hex_char;
			L30_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_22;
--sw  R24 [] 
--dw  R24 [] 
--sc  R24 [] 
--lc  R24 [] 
	component route_23 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne992 : in hex_char;
			ne992_command : out routeCommands := RELEASE;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			J40_state : in hex_char;
			J40_command : out routeCommands := RELEASE;
			L31_state : in hex_char;
			L31_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_23;
--sw  R25 [] 
--dw  R25 [] 
--sc  R25 [] 
--lc  R25 [] 
	component route_24 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			J43_state : in hex_char;
			J43_command : out routeCommands := RELEASE;
			X53_state : in hex_char;
			X53_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_24;
--sw  R26 ['D09'] 
--dw  R26 [] 
--sc  R26 [] 
--lc  R26 [] 
	component route_25 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne912 : in hex_char;
			ne912_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			J45_state : in hex_char;
			J45_command : out routeCommands := RELEASE;
			J43_state : in hex_char;
			J43_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_25;
--sw  R27 ['D23'] 
--dw  R27 [] 
--sc  R27 [] 
--lc  R27 [] 
	component route_26 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne132 : in hex_char;
			ne132_command : out routeCommands := RELEASE;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			J46_state : in hex_char;
			J46_command : out routeCommands := RELEASE;
			L29_state : in hex_char;
			L29_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_26;
--sw  R28 ['D09', 'D20'] 
--dw  R28 [] 
--sc  R28 [] 
--lc  R28 [] 
	component route_27 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne132 : in hex_char;
			ne132_command : out routeCommands := RELEASE;
			track_ne912 : in hex_char;
			ne912_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D20_state : in hex_char;
			D20_command : out routeCommands := RELEASE;
			J47_state : in hex_char;
			J47_command : out routeCommands := RELEASE;
			J45_state : in hex_char;
			J45_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_27;
--sw  R29 [] 
--dw  R29 [] 
--sc  R29 [] 
--lc  R29 [] 
	component route_28 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			track_ne102 : in hex_char;
			ne102_command : out routeCommands := RELEASE;
			J48_state : in hex_char;
			J48_command : out routeCommands := RELEASE;
			T11_state : in hex_char;
			T11_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_28;
--sw  R30 ['D05'] 
--dw  R30 [] 
--sc  R30 [] 
--lc  R30 ['Lc01'] 
	component route_29 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			X50_state : in hex_char;
			X50_command : out routeCommands := RELEASE;
			S55_state : in hex_char;
			S55_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_29;
--sw  R31 ['Sw04', 'Sw03'] 
--dw  R31 [] 
--sc  R31 [] 
--lc  R31 ['Lc01'] 
	component route_30 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			track_ne996 : in hex_char;
			ne996_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			X51_state : in hex_char;
			X51_command : out routeCommands := RELEASE;
			S129_state : in hex_char;
			S129_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_30;
--sw  R32 ['D09'] 
--dw  R32 [] 
--sc  R32 [] 
--lc  R32 ['Lc04'] 
	component route_31 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			Lc04_state : in hex_char;
			Lc04_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			X52_state : in hex_char;
			X52_command : out routeCommands := RELEASE;
			S59_state : in hex_char;
			S59_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_31;
--sw  R33 ['Sw01', 'Sw05'] 
--dw  R33 [] 
--sc  R33 [] 
--lc  R33 ['Lc04'] 
	component route_32 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			track_ne992 : in hex_char;
			ne992_command : out routeCommands := RELEASE;
			Lc04_state : in hex_char;
			Lc04_command : out routeCommands := RELEASE;
			Sw01_state : in hex_char;
			Sw01_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			X53_state : in hex_char;
			X53_command : out routeCommands := RELEASE;
			S120_state : in hex_char;
			S120_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_32;
--sw  R34 ['D05'] 
--dw  R34 [] 
--sc  R34 [] 
--lc  R34 ['Lc01'] 
	component route_33 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne63 : in hex_char;
			ne63_command : out routeCommands := RELEASE;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			C54_state : in hex_char;
			C54_command : out routeCommands := RELEASE;
			X51_state : in hex_char;
			X51_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_33;
--sw  R35 ['D08', 'D05'] 
--dw  R35 [] 
--sc  R35 [] 
--lc  R35 [] 
	component route_34 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			track_ne61 : in hex_char;
			ne61_command : out routeCommands := RELEASE;
			D08_state : in hex_char;
			D08_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			S55_state : in hex_char;
			S55_command : out routeCommands := RELEASE;
			S78_state : in hex_char;
			S78_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_34;
--sw  R36 ['D05', 'D18'] 
--dw  R36 [] 
--sc  R36 [] 
--lc  R36 [] 
	component route_35 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			track_ne63 : in hex_char;
			ne63_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			D18_state : in hex_char;
			D18_command : out routeCommands := RELEASE;
			S55_state : in hex_char;
			S55_command : out routeCommands := RELEASE;
			S95_state : in hex_char;
			S95_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_35;
--sw  R37 ['D09', 'D20', 'D21'] 
--dw  R37 [] 
--sc  R37 [] 
--lc  R37 [] 
	component route_36 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			track_ne912 : in hex_char;
			ne912_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D20_state : in hex_char;
			D20_command : out routeCommands := RELEASE;
			D21_state : in hex_char;
			D21_command : out routeCommands := RELEASE;
			S59_state : in hex_char;
			S59_command : out routeCommands := RELEASE;
			S110_state : in hex_char;
			S110_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_36;
--sw  R38 ['D10', 'D09'] 
--dw  R38 [] 
--sc  R38 [] 
--lc  R38 [] 
	component route_37 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			track_ne910 : in hex_char;
			ne910_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			S59_state : in hex_char;
			S59_command : out routeCommands := RELEASE;
			S81_state : in hex_char;
			S81_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_37;
--sw  R39 ['D01', 'D03'] 
--dw  R39 [] 
--sc  R39 [] 
--lc  R39 [] 
	component route_38 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne991 : in hex_char;
			ne991_command : out routeCommands := RELEASE;
			track_ne288 : in hex_char;
			ne288_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			D03_state : in hex_char;
			D03_command : out routeCommands := RELEASE;
			S64_state : in hex_char;
			S64_command : out routeCommands := RELEASE;
			S69_state : in hex_char;
			S69_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_38;
--sw  R40 ['D01', 'D14'] 
--dw  R40 [] 
--sc  R40 [] 
--lc  R40 [] 
	component route_39 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne991 : in hex_char;
			ne991_command : out routeCommands := RELEASE;
			track_ne290 : in hex_char;
			ne290_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			D14_state : in hex_char;
			D14_command : out routeCommands := RELEASE;
			S64_state : in hex_char;
			S64_command : out routeCommands := RELEASE;
			S86_state : in hex_char;
			S86_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_39;
--sw  R41 ['D01', 'D03'] 
--dw  R41 [] 
--sc  R41 [] 
--lc  R41 [] 
	component route_40 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne295 : in hex_char;
			ne295_command : out routeCommands := RELEASE;
			track_ne288 : in hex_char;
			ne288_command : out routeCommands := RELEASE;
			track_ne991 : in hex_char;
			ne991_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			D03_state : in hex_char;
			D03_command : out routeCommands := RELEASE;
			C67_state : in hex_char;
			C67_command : out routeCommands := RELEASE;
			T01_state : in hex_char;
			T01_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_40;
--sw  R42 ['D04', 'Sw03', 'Sw02'] 
--dw  R42 [] 
--sc  R42 [] 
--lc  R42 [] 
	component route_41 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			track_ne384 : in hex_char;
			ne384_command : out routeCommands := RELEASE;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			Sw02_state : in hex_char;
			Sw02_command : out routeCommands := RELEASE;
			B68_state : in hex_char;
			B68_command : out routeCommands := RELEASE;
			S126_state : in hex_char;
			S126_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_41;
--sw  R43 ['D03', 'D04'] 
--dw  R43 [] 
--sc  R43 [] 
--lc  R43 [] 
	component route_42 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne288 : in hex_char;
			ne288_command : out routeCommands := RELEASE;
			track_ne295 : in hex_char;
			ne295_command : out routeCommands := RELEASE;
			D03_state : in hex_char;
			D03_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			S69_state : in hex_char;
			S69_command : out routeCommands := RELEASE;
			C70_state : in hex_char;
			C70_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_42;
--sw  R44 ['D03', 'D04', 'Sw02'] 
--dw  R44 [] 
--sc  R44 [] 
--lc  R44 [] 
	component route_43 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne288 : in hex_char;
			ne288_command : out routeCommands := RELEASE;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			D03_state : in hex_char;
			D03_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			Sw02_state : in hex_char;
			Sw02_command : out routeCommands := RELEASE;
			S69_state : in hex_char;
			S69_command : out routeCommands := RELEASE;
			B68_state : in hex_char;
			B68_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_43;
--sw  R45 ['D04', 'Sw03'] 
--dw  R45 [] 
--sc  R45 [] 
--lc  R45 [] 
	component route_44 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne295 : in hex_char;
			ne295_command : out routeCommands := RELEASE;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			C70_state : in hex_char;
			C70_command : out routeCommands := RELEASE;
			S126_state : in hex_char;
			S126_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_44;
--sw  R46 ['D01', 'D03', 'D04'] 
--dw  R46 [] 
--sc  R46 [] 
--lc  R46 [] 
	component route_45 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			track_ne295 : in hex_char;
			ne295_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			D03_state : in hex_char;
			D03_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			S71_state : in hex_char;
			S71_command : out routeCommands := RELEASE;
			C67_state : in hex_char;
			C67_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_45;
--sw  R47 ['D04', 'Sw02'] 
--dw  R47 [] 
--sc  R47 [] 
--lc  R47 [] 
	component route_46 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			track_ne384 : in hex_char;
			ne384_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			Sw02_state : in hex_char;
			Sw02_command : out routeCommands := RELEASE;
			S71_state : in hex_char;
			S71_command : out routeCommands := RELEASE;
			S84_state : in hex_char;
			S84_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_46;
--sw  R48 ['D07', 'Sw05'] 
--dw  R48 [] 
--sc  R48 [] 
--lc  R48 [] 
	component route_47 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne404 : in hex_char;
			ne404_command : out routeCommands := RELEASE;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			C73_state : in hex_char;
			C73_command : out routeCommands := RELEASE;
			S123_state : in hex_char;
			S123_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_47;
--sw  R49 ['D08', 'D05', 'D07'] 
--dw  R49 [] 
--sc  R49 [] 
--lc  R49 [] 
	component route_48 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			track_ne404 : in hex_char;
			ne404_command : out routeCommands := RELEASE;
			D08_state : in hex_char;
			D08_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			S74_state : in hex_char;
			S74_command : out routeCommands := RELEASE;
			C76_state : in hex_char;
			C76_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_48;
--sw  R50 ['D07', 'D16'] 
--dw  R50 [] 
--sc  R50 [] 
--lc  R50 [] 
	component route_49 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			track_ne407 : in hex_char;
			ne407_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			D16_state : in hex_char;
			D16_command : out routeCommands := RELEASE;
			S74_state : in hex_char;
			S74_command : out routeCommands := RELEASE;
			S93_state : in hex_char;
			S93_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_49;
--sw  R51 ['D08', 'D05'] 
--dw  R51 [] 
--sc  R51 [] 
--lc  R51 ['Lc01'] 
	component route_50 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne404 : in hex_char;
			ne404_command : out routeCommands := RELEASE;
			track_ne61 : in hex_char;
			ne61_command : out routeCommands := RELEASE;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			D08_state : in hex_char;
			D08_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			C76_state : in hex_char;
			C76_command : out routeCommands := RELEASE;
			X51_state : in hex_char;
			X51_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_50;
--sw  R52 ['D07', 'Sw05', 'D16'] 
--dw  R52 [] 
--sc  R52 [] 
--lc  R52 [] 
	component route_51 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne123 : in hex_char;
			ne123_command : out routeCommands := RELEASE;
			track_ne407 : in hex_char;
			ne407_command : out routeCommands := RELEASE;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			D16_state : in hex_char;
			D16_command : out routeCommands := RELEASE;
			B77_state : in hex_char;
			B77_command : out routeCommands := RELEASE;
			S123_state : in hex_char;
			S123_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_51;
--sw  R53 ['D08', 'D07'] 
--dw  R53 [] 
--sc  R53 [] 
--lc  R53 [] 
	component route_52 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne61 : in hex_char;
			ne61_command : out routeCommands := RELEASE;
			track_ne404 : in hex_char;
			ne404_command : out routeCommands := RELEASE;
			D08_state : in hex_char;
			D08_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			S78_state : in hex_char;
			S78_command : out routeCommands := RELEASE;
			C73_state : in hex_char;
			C73_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_52;
--sw  R54 ['D08', 'D07', 'D16'] 
--dw  R54 [] 
--sc  R54 [] 
--lc  R54 [] 
	component route_53 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne61 : in hex_char;
			ne61_command : out routeCommands := RELEASE;
			track_ne123 : in hex_char;
			ne123_command : out routeCommands := RELEASE;
			D08_state : in hex_char;
			D08_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			D16_state : in hex_char;
			D16_command : out routeCommands := RELEASE;
			S78_state : in hex_char;
			S78_command : out routeCommands := RELEASE;
			B77_state : in hex_char;
			B77_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_53;
--sw  R55 ['D10', 'D09'] 
--dw  R55 [] 
--sc  R55 [] 
--lc  R55 [] 
	component route_54 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne130 : in hex_char;
			ne130_command : out routeCommands := RELEASE;
			track_ne910 : in hex_char;
			ne910_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			C79_state : in hex_char;
			C79_command : out routeCommands := RELEASE;
			J43_state : in hex_char;
			J43_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_54;
--sw  R56 ['D23', 'D24'] 
--dw  R56 [] 
--sc  R56 [] 
--lc  R56 [] 
	component route_55 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne135 : in hex_char;
			ne135_command : out routeCommands := RELEASE;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			D24_state : in hex_char;
			D24_command : out routeCommands := RELEASE;
			B80_state : in hex_char;
			B80_command : out routeCommands := RELEASE;
			S104_state : in hex_char;
			S104_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_55;
--sw  R57 ['D10', 'D23'] 
--dw  R57 [] 
--sc  R57 [] 
--lc  R57 [] 
	component route_56 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne910 : in hex_char;
			ne910_command : out routeCommands := RELEASE;
			track_ne130 : in hex_char;
			ne130_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			S81_state : in hex_char;
			S81_command : out routeCommands := RELEASE;
			S107_state : in hex_char;
			S107_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_56;
--sw  R58 ['D10', 'D24'] 
--dw  R58 [] 
--sc  R58 [] 
--lc  R58 [] 
	component route_57 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne910 : in hex_char;
			ne910_command : out routeCommands := RELEASE;
			track_ne135 : in hex_char;
			ne135_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D24_state : in hex_char;
			D24_command : out routeCommands := RELEASE;
			S81_state : in hex_char;
			S81_command : out routeCommands := RELEASE;
			B80_state : in hex_char;
			B80_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_57;
--sw  R59 ['Sw02'] 
--dw  R59 [] 
--sc  R59 [] 
--lc  R59 [] 
	component route_58 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne384 : in hex_char;
			ne384_command : out routeCommands := RELEASE;
			track_ne104 : in hex_char;
			ne104_command : out routeCommands := RELEASE;
			Sw02_state : in hex_char;
			Sw02_command : out routeCommands := RELEASE;
			S84_state : in hex_char;
			S84_command : out routeCommands := RELEASE;
			T13_state : in hex_char;
			T13_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_58;
--sw  R60 ['D01', 'D03', 'Sw02'] 
--dw  R60 [] 
--sc  R60 [] 
--lc  R60 [] 
	component route_59 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne384 : in hex_char;
			ne384_command : out routeCommands := RELEASE;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			track_ne288 : in hex_char;
			ne288_command : out routeCommands := RELEASE;
			track_ne991 : in hex_char;
			ne991_command : out routeCommands := RELEASE;
			D01_state : in hex_char;
			D01_command : out routeCommands := RELEASE;
			D03_state : in hex_char;
			D03_command : out routeCommands := RELEASE;
			Sw02_state : in hex_char;
			Sw02_command : out routeCommands := RELEASE;
			S84_state : in hex_char;
			S84_command : out routeCommands := RELEASE;
			T01_state : in hex_char;
			T01_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_59;
--sw  R61 ['D14', 'Sw04'] 
--dw  R61 [] 
--sc  R61 [] 
--lc  R61 [] 
	component route_60 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne290 : in hex_char;
			ne290_command : out routeCommands := RELEASE;
			track_ne292 : in hex_char;
			ne292_command : out routeCommands := RELEASE;
			D14_state : in hex_char;
			D14_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			S86_state : in hex_char;
			S86_command : out routeCommands := RELEASE;
			J36_state : in hex_char;
			J36_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_60;
--sw  R62 ['D14', 'D15'] 
--dw  R62 [] 
--sc  R62 [] 
--lc  R62 [] 
	component route_61 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne290 : in hex_char;
			ne290_command : out routeCommands := RELEASE;
			track_ne111 : in hex_char;
			ne111_command : out routeCommands := RELEASE;
			track_ne377 : in hex_char;
			ne377_command : out routeCommands := RELEASE;
			D14_state : in hex_char;
			D14_command : out routeCommands := RELEASE;
			D15_state : in hex_char;
			D15_command : out routeCommands := RELEASE;
			S86_state : in hex_char;
			S86_command : out routeCommands := RELEASE;
			T03_state : in hex_char;
			T03_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_61;
--sw  R63 ['D16'] 
--dw  R63 [] 
--sc  R63 [] 
--lc  R63 [] 
	component route_62 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne407 : in hex_char;
			ne407_command : out routeCommands := RELEASE;
			track_ne122 : in hex_char;
			ne122_command : out routeCommands := RELEASE;
			D16_state : in hex_char;
			D16_command : out routeCommands := RELEASE;
			S93_state : in hex_char;
			S93_command : out routeCommands := RELEASE;
			T17_state : in hex_char;
			T17_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_62;
--sw  R64 ['D08', 'D05', 'D16'] 
--dw  R64 [] 
--sc  R64 [] 
--lc  R64 ['Lc01'] 
	component route_63 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne407 : in hex_char;
			ne407_command : out routeCommands := RELEASE;
			track_ne123 : in hex_char;
			ne123_command : out routeCommands := RELEASE;
			track_ne61 : in hex_char;
			ne61_command : out routeCommands := RELEASE;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			D08_state : in hex_char;
			D08_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			D16_state : in hex_char;
			D16_command : out routeCommands := RELEASE;
			S93_state : in hex_char;
			S93_command : out routeCommands := RELEASE;
			X51_state : in hex_char;
			X51_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_63;
--sw  R65 ['D05', 'D18'] 
--dw  R65 [] 
--sc  R65 [] 
--lc  R65 [] 
	component route_64 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne65 : in hex_char;
			ne65_command : out routeCommands := RELEASE;
			track_ne63 : in hex_char;
			ne63_command : out routeCommands := RELEASE;
			D05_state : in hex_char;
			D05_command : out routeCommands := RELEASE;
			D18_state : in hex_char;
			D18_command : out routeCommands := RELEASE;
			C94_state : in hex_char;
			C94_command : out routeCommands := RELEASE;
			C54_state : in hex_char;
			C54_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_64;
--sw  R66 ['D18', 'Sw01'] 
--dw  R66 [] 
--sc  R66 [] 
--lc  R66 [] 
	component route_65 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne63 : in hex_char;
			ne63_command : out routeCommands := RELEASE;
			track_ne65 : in hex_char;
			ne65_command : out routeCommands := RELEASE;
			D18_state : in hex_char;
			D18_command : out routeCommands := RELEASE;
			Sw01_state : in hex_char;
			Sw01_command : out routeCommands := RELEASE;
			S95_state : in hex_char;
			S95_command : out routeCommands := RELEASE;
			C119_state : in hex_char;
			C119_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_65;
--sw  R67 ['D18', 'D19'] 
--dw  R67 [] 
--sc  R67 [] 
--lc  R67 [] 
	component route_66 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne63 : in hex_char;
			ne63_command : out routeCommands := RELEASE;
			track_ne124 : in hex_char;
			ne124_command : out routeCommands := RELEASE;
			track_ne421 : in hex_char;
			ne421_command : out routeCommands := RELEASE;
			D18_state : in hex_char;
			D18_command : out routeCommands := RELEASE;
			D19_state : in hex_char;
			D19_command : out routeCommands := RELEASE;
			S95_state : in hex_char;
			S95_command : out routeCommands := RELEASE;
			T05_state : in hex_char;
			T05_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_66;
--sw  R68 ['D20', 'D23'] 
--dw  R68 [] 
--sc  R68 [] 
--lc  R68 [] 
	component route_67 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			track_ne132 : in hex_char;
			ne132_command : out routeCommands := RELEASE;
			D20_state : in hex_char;
			D20_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			S101_state : in hex_char;
			S101_command : out routeCommands := RELEASE;
			J47_state : in hex_char;
			J47_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_67;
--sw  R69 ['D10', 'D09', 'D23', 'D24'] 
--dw  R69 ['D12'] 
--sc  R69 [] 
--lc  R69 [] 
	component route_68 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			track_ne129 : in hex_char;
			ne129_command : out routeCommands := RELEASE;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			D24_state : in hex_char;
			D24_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			S101_state : in hex_char;
			S101_command : out routeCommands := RELEASE;
			S117_state : in hex_char;
			S117_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_68;
--sw  R70 ['D10', 'D09', 'D23'] 
--dw  R70 ['D12'] 
--sc  R70 [] 
--lc  R70 [] 
	component route_69 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			track_ne129 : in hex_char;
			ne129_command : out routeCommands := RELEASE;
			track_ne130 : in hex_char;
			ne130_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			S101_state : in hex_char;
			S101_command : out routeCommands := RELEASE;
			C79_state : in hex_char;
			C79_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_69;
--sw  R71 ['D23'] 
--dw  R71 ['D12'] 
--sc  R71 [] 
--lc  R71 [] 
	component route_70 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			track_ne129 : in hex_char;
			ne129_command : out routeCommands := RELEASE;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			S104_state : in hex_char;
			S104_command : out routeCommands := RELEASE;
			L29_state : in hex_char;
			L29_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_70;
--sw  R72 [] 
--dw  R72 ['D12'] 
--sc  R72 [] 
--lc  R72 [] 
	component route_71 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			track_ne450 : in hex_char;
			ne450_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			S104_state : in hex_char;
			S104_command : out routeCommands := RELEASE;
			T07_state : in hex_char;
			T07_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_71;
--sw  R73 ['D23'] 
--dw  R73 ['D12'] 
--sc  R73 [] 
--lc  R73 [] 
	component route_72 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne130 : in hex_char;
			ne130_command : out routeCommands := RELEASE;
			track_ne129 : in hex_char;
			ne129_command : out routeCommands := RELEASE;
			track_ne114 : in hex_char;
			ne114_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			S107_state : in hex_char;
			S107_command : out routeCommands := RELEASE;
			L29_state : in hex_char;
			L29_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_72;
--sw  R74 [] 
--dw  R74 ['D12'] 
--sc  R74 [] 
--lc  R74 [] 
	component route_73 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne130 : in hex_char;
			ne130_command : out routeCommands := RELEASE;
			track_ne450 : in hex_char;
			ne450_command : out routeCommands := RELEASE;
			D12_state : in hex_char;
			D12_command : out routeCommands := RELEASE;
			S107_state : in hex_char;
			S107_command : out routeCommands := RELEASE;
			T07_state : in hex_char;
			T07_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_73;
--sw  R75 ['D20', 'D21'] 
--dw  R75 [] 
--sc  R75 [] 
--lc  R75 [] 
	component route_74 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne912 : in hex_char;
			ne912_command : out routeCommands := RELEASE;
			track_ne131 : in hex_char;
			ne131_command : out routeCommands := RELEASE;
			track_ne465 : in hex_char;
			ne465_command : out routeCommands := RELEASE;
			D20_state : in hex_char;
			D20_command : out routeCommands := RELEASE;
			D21_state : in hex_char;
			D21_command : out routeCommands := RELEASE;
			S110_state : in hex_char;
			S110_command : out routeCommands := RELEASE;
			T09_state : in hex_char;
			T09_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_74;
--sw  R76 ['D20', 'D23'] 
--dw  R76 [] 
--sc  R76 [] 
--lc  R76 [] 
	component route_75 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne912 : in hex_char;
			ne912_command : out routeCommands := RELEASE;
			track_ne132 : in hex_char;
			ne132_command : out routeCommands := RELEASE;
			D20_state : in hex_char;
			D20_command : out routeCommands := RELEASE;
			D23_state : in hex_char;
			D23_command : out routeCommands := RELEASE;
			S110_state : in hex_char;
			S110_command : out routeCommands := RELEASE;
			J46_state : in hex_char;
			J46_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_75;
--sw  R77 ['D10', 'D09', 'D24'] 
--dw  R77 [] 
--sc  R77 [] 
--lc  R77 [] 
	component route_76 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			track_ne135 : in hex_char;
			ne135_command : out routeCommands := RELEASE;
			track_ne910 : in hex_char;
			ne910_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			D10_state : in hex_char;
			D10_command : out routeCommands := RELEASE;
			D09_state : in hex_char;
			D09_command : out routeCommands := RELEASE;
			D24_state : in hex_char;
			D24_command : out routeCommands := RELEASE;
			S117_state : in hex_char;
			S117_command : out routeCommands := RELEASE;
			J43_state : in hex_char;
			J43_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_76;
--sw  R78 ['D24'] 
--dw  R78 [] 
--sc  R78 [] 
--lc  R78 [] 
	component route_77 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne127 : in hex_char;
			ne127_command : out routeCommands := RELEASE;
			track_ne134 : in hex_char;
			ne134_command : out routeCommands := RELEASE;
			D24_state : in hex_char;
			D24_command : out routeCommands := RELEASE;
			S117_state : in hex_char;
			S117_command : out routeCommands := RELEASE;
			T23_state : in hex_char;
			T23_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_77;
--sw  R79 ['Sw01'] 
--dw  R79 [] 
--sc  R79 [] 
--lc  R79 [] 
	component route_78 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne65 : in hex_char;
			ne65_command : out routeCommands := RELEASE;
			track_ne992 : in hex_char;
			ne992_command : out routeCommands := RELEASE;
			Sw01_state : in hex_char;
			Sw01_command : out routeCommands := RELEASE;
			C119_state : in hex_char;
			C119_command : out routeCommands := RELEASE;
			J40_state : in hex_char;
			J40_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_78;
--sw  R80 ['D18', 'Sw01'] 
--dw  R80 [] 
--sc  R80 [] 
--lc  R80 [] 
	component route_79 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne992 : in hex_char;
			ne992_command : out routeCommands := RELEASE;
			track_ne65 : in hex_char;
			ne65_command : out routeCommands := RELEASE;
			D18_state : in hex_char;
			D18_command : out routeCommands := RELEASE;
			Sw01_state : in hex_char;
			Sw01_command : out routeCommands := RELEASE;
			S120_state : in hex_char;
			S120_command : out routeCommands := RELEASE;
			C94_state : in hex_char;
			C94_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_79;
--sw  R81 ['Sw01', 'D07', 'Sw05'] 
--dw  R81 [] 
--sc  R81 [] 
--lc  R81 [] 
	component route_80 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne992 : in hex_char;
			ne992_command : out routeCommands := RELEASE;
			track_ne994 : in hex_char;
			ne994_command : out routeCommands := RELEASE;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			Sw01_state : in hex_char;
			Sw01_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			S120_state : in hex_char;
			S120_command : out routeCommands := RELEASE;
			S74_state : in hex_char;
			S74_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_80;
--sw  R82 ['D07', 'Sw05'] 
--dw  R82 [] 
--sc  R82 [] 
--lc  R82 [] 
	component route_81 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne993 : in hex_char;
			ne993_command : out routeCommands := RELEASE;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			D07_state : in hex_char;
			D07_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			C122_state : in hex_char;
			C122_command : out routeCommands := RELEASE;
			S74_state : in hex_char;
			S74_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_81;
--sw  R83 ['Sw05'] 
--dw  R83 [] 
--sc  R83 [] 
--lc  R83 [] 
	component route_82 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			track_ne993 : in hex_char;
			ne993_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			S123_state : in hex_char;
			S123_command : out routeCommands := RELEASE;
			T25_state : in hex_char;
			T25_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_82;
--sw  R84 ['Sw01', 'Sw05'] 
--dw  R84 [] 
--sc  R84 [] 
--lc  R84 [] 
	component route_83 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne400 : in hex_char;
			ne400_command : out routeCommands := RELEASE;
			track_ne994 : in hex_char;
			ne994_command : out routeCommands := RELEASE;
			track_ne992 : in hex_char;
			ne992_command : out routeCommands := RELEASE;
			Sw01_state : in hex_char;
			Sw01_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			S123_state : in hex_char;
			S123_command : out routeCommands := RELEASE;
			J40_state : in hex_char;
			J40_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_83;
--sw  R85 ['D04', 'Sw03'] 
--dw  R85 [] 
--sc  R85 [] 
--lc  R85 [] 
	component route_84 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne995 : in hex_char;
			ne995_command : out routeCommands := RELEASE;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			C125_state : in hex_char;
			C125_command : out routeCommands := RELEASE;
			S71_state : in hex_char;
			S71_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_84;
--sw  R86 ['Sw03'] 
--dw  R86 [] 
--sc  R86 [] 
--lc  R86 [] 
	component route_85 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			track_ne995 : in hex_char;
			ne995_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			S126_state : in hex_char;
			S126_command : out routeCommands := RELEASE;
			T27_state : in hex_char;
			T27_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_85;
--sw  R87 ['Sw04', 'Sw03'] 
--dw  R87 [] 
--sc  R87 [] 
--lc  R87 [] 
	component route_86 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			track_ne997 : in hex_char;
			ne997_command : out routeCommands := RELEASE;
			track_ne996 : in hex_char;
			ne996_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			S126_state : in hex_char;
			S126_command : out routeCommands := RELEASE;
			J38_state : in hex_char;
			J38_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_86;
--sw  R88 ['D14', 'Sw04'] 
--dw  R88 [] 
--sc  R88 [] 
--lc  R88 [] 
	component route_87 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne996 : in hex_char;
			ne996_command : out routeCommands := RELEASE;
			track_ne292 : in hex_char;
			ne292_command : out routeCommands := RELEASE;
			D14_state : in hex_char;
			D14_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			S129_state : in hex_char;
			S129_command : out routeCommands := RELEASE;
			J37_state : in hex_char;
			J37_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_87;
--sw  R89 ['Sw04', 'D04', 'Sw03'] 
--dw  R89 [] 
--sc  R89 [] 
--lc  R89 [] 
	component route_88 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne996 : in hex_char;
			ne996_command : out routeCommands := RELEASE;
			track_ne997 : in hex_char;
			ne997_command : out routeCommands := RELEASE;
			track_ne297 : in hex_char;
			ne297_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			D04_state : in hex_char;
			D04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			S129_state : in hex_char;
			S129_command : out routeCommands := RELEASE;
			S71_state : in hex_char;
			S71_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_88;
	signal state_Lc01 , state_Lc04 : hex_char;
	signal state_D01 , state_D08 , state_D05 , state_D18 , state_Sw01 , state_D10 , state_D09 , state_D20 , state_D23 , state_D03 , state_D14 , state_Sw04 , state_D04 , state_Sw03 , state_D15 , state_Sw02 , state_D07 , state_Sw05 , state_D16 , state_D19 , state_D21 , state_D24 : hex_char;
	signal state_D12 : hex_char;
	signal state_T01 , state_T02 , state_S64 , state_S78 , state_C54 , state_S95 , state_C94 , state_C119 , state_S81 , state_J45 , state_S110 , state_L29 , state_J48 , state_S101 , state_S69 , state_J35 , state_S86 , state_J36 , state_J37 , state_C67 , state_C70 , state_S71 , state_S126 , state_T03 , state_T04 , state_S84 , state_S74 , state_S123 , state_C73 , state_C76 , state_S93 , state_T05 , state_T06 , state_T07 , state_T08 , state_T09 , state_T10 , state_L30 , state_X50 , state_X51 , state_S55 , state_L31 , state_X52 , state_X53 , state_J43 , state_S59 , state_T11 , state_T12 , state_T13 , state_T14 , state_B68 , state_T15 , state_T16 , state_T17 , state_T18 , state_B77 , state_T19 , state_T20 , state_S104 , state_S117 , state_C79 , state_S107 , state_J46 , state_J47 , state_T21 , state_T22 , state_T23 , state_T24 , state_B80 , state_J40 , state_S120 , state_T25 , state_C122 , state_T27 , state_C125 , state_J38 , state_S129 : hex_char;
	signal cmd_R1_ne991 , cmd_R2_ne377 , cmd_R2_ne111 , cmd_R2_ne290 , cmd_R3_ne377 , cmd_R3_ne113 , cmd_R4_ne421 , cmd_R4_ne124 , cmd_R4_ne63 , cmd_R5_ne421 , cmd_R5_ne126 , cmd_R6_ne450 , cmd_R6_ne127 , cmd_R7_ne450 , cmd_R7_ne130 , cmd_R8_ne465 , cmd_R8_ne131 , cmd_R8_ne912 , cmd_R9_ne465 , cmd_R9_ne133 , cmd_R10_ne102 , cmd_R10_ne114 , cmd_R11_ne104 , cmd_R11_ne384 , cmd_R11_ne297 , cmd_R12_ne113 , cmd_R12_ne377 , cmd_R13_ne122 , cmd_R13_ne407 , cmd_R13_ne400 , cmd_R14_ne126 , cmd_R14_ne421 , cmd_R15_ne133 , cmd_R15_ne465 , cmd_R16_ne134 , cmd_R16_ne127 , cmd_R17_ne114 , cmd_R18_ne98 , cmd_R19_ne100 , cmd_R20_ne290 , cmd_R20_ne991 , cmd_R21_ne292 , cmd_R21_ne996 , cmd_R22_ne292 , cmd_R22_ne290 , cmd_R23_ne996 , cmd_R23_ne98 , cmd_R24_ne992 , cmd_R24_ne100 , cmd_R25_ne101 , cmd_R25_ne100 , cmd_R26_ne912 , cmd_R26_ne101 , cmd_R27_ne132 , cmd_R27_ne114 , cmd_R28_ne132 , cmd_R28_ne912 , cmd_R29_ne114 , cmd_R29_ne102 , cmd_R30_ne98 , cmd_R30_ne99 , cmd_R31_ne98 , cmd_R31_ne996 , cmd_R32_ne100 , cmd_R32_ne101 , cmd_R33_ne100 , cmd_R33_ne992 , cmd_R34_ne63 , cmd_R34_ne99 , cmd_R34_ne98 , cmd_R35_ne99 , cmd_R35_ne61 , cmd_R36_ne99 , cmd_R36_ne63 , cmd_R37_ne101 , cmd_R37_ne912 , cmd_R38_ne101 , cmd_R38_ne910 , cmd_R39_ne991 , cmd_R39_ne288 , cmd_R40_ne991 , cmd_R40_ne290 , cmd_R41_ne295 , cmd_R41_ne288 , cmd_R41_ne991 , cmd_R42_ne110 , cmd_R42_ne384 , cmd_R42_ne297 , cmd_R43_ne288 , cmd_R43_ne295 , cmd_R44_ne288 , cmd_R44_ne110 , cmd_R45_ne295 , cmd_R45_ne297 , cmd_R46_ne297 , cmd_R46_ne295 , cmd_R47_ne297 , cmd_R47_ne384 , cmd_R48_ne404 , cmd_R48_ne400 , cmd_R49_ne400 , cmd_R49_ne404 , cmd_R50_ne400 , cmd_R50_ne407 , cmd_R51_ne404 , cmd_R51_ne61 , cmd_R51_ne99 , cmd_R51_ne98 , cmd_R52_ne123 , cmd_R52_ne407 , cmd_R52_ne400 , cmd_R53_ne61 , cmd_R53_ne404 , cmd_R54_ne61 , cmd_R54_ne123 , cmd_R55_ne130 , cmd_R55_ne910 , cmd_R55_ne101 , cmd_R56_ne135 , cmd_R56_ne127 , cmd_R57_ne910 , cmd_R57_ne130 , cmd_R58_ne910 , cmd_R58_ne135 , cmd_R59_ne384 , cmd_R59_ne104 , cmd_R60_ne384 , cmd_R60_ne110 , cmd_R60_ne288 , cmd_R60_ne991 , cmd_R61_ne290 , cmd_R61_ne292 , cmd_R62_ne290 , cmd_R62_ne111 , cmd_R62_ne377 , cmd_R63_ne407 , cmd_R63_ne122 , cmd_R64_ne407 , cmd_R64_ne123 , cmd_R64_ne61 , cmd_R64_ne99 , cmd_R64_ne98 , cmd_R65_ne65 , cmd_R65_ne63 , cmd_R66_ne63 , cmd_R66_ne65 , cmd_R67_ne63 , cmd_R67_ne124 , cmd_R67_ne421 , cmd_R68_ne114 , cmd_R68_ne132 , cmd_R69_ne114 , cmd_R69_ne129 , cmd_R69_ne127 , cmd_R70_ne114 , cmd_R70_ne129 , cmd_R70_ne130 , cmd_R71_ne127 , cmd_R71_ne129 , cmd_R71_ne114 , cmd_R72_ne127 , cmd_R72_ne450 , cmd_R73_ne130 , cmd_R73_ne129 , cmd_R73_ne114 , cmd_R74_ne130 , cmd_R74_ne450 , cmd_R75_ne912 , cmd_R75_ne131 , cmd_R75_ne465 , cmd_R76_ne912 , cmd_R76_ne132 , cmd_R77_ne127 , cmd_R77_ne135 , cmd_R77_ne910 , cmd_R77_ne101 , cmd_R78_ne127 , cmd_R78_ne134 , cmd_R79_ne65 , cmd_R79_ne992 , cmd_R80_ne992 , cmd_R80_ne65 , cmd_R81_ne992 , cmd_R81_ne994 , cmd_R81_ne400 , cmd_R82_ne993 , cmd_R82_ne400 , cmd_R83_ne400 , cmd_R83_ne993 , cmd_R84_ne400 , cmd_R84_ne994 , cmd_R84_ne992 , cmd_R85_ne995 , cmd_R85_ne297 , cmd_R86_ne297 , cmd_R86_ne995 , cmd_R87_ne297 , cmd_R87_ne997 , cmd_R87_ne996 , cmd_R88_ne996 , cmd_R88_ne292 , cmd_R89_ne996 , cmd_R89_ne997 , cmd_R89_ne297 : routeCommands := RELEASE;
	signal state_ne991 , state_ne61 , state_ne63 , state_ne65 , state_ne910 , state_ne912 , state_ne114 , state_ne288 , state_ne290 , state_ne292 , state_ne295 , state_ne297 , state_ne377 , state_ne384 , state_ne400 , state_ne404 , state_ne407 , state_ne421 , state_ne450 , state_ne465 , state_ne98 , state_ne99 , state_ne100 , state_ne101 , state_ne102 , state_ne104 , state_ne110 , state_ne111 , state_ne113 , state_ne122 , state_ne123 , state_ne124 , state_ne126 , state_ne127 , state_ne129 , state_ne130 , state_ne131 , state_ne132 , state_ne133 , state_ne134 , state_ne135 , state_ne992 , state_ne993 , state_ne994 , state_ne995 , state_ne996 , state_ne997 : hex_char;
	signal cmd_R30_Lc01 , cmd_R31_Lc01 , cmd_R34_Lc01 , cmd_R51_Lc01 , cmd_R64_Lc01 , cmd_R32_Lc04 , cmd_R33_Lc04 : routeCommands := RELEASE;
	signal cmd_R20_D01 , cmd_R39_D01 , cmd_R40_D01 , cmd_R41_D01 , cmd_R60_D01 , cmd_R1_D01 , cmd_R22_D01 , cmd_R46_D01 , cmd_R2_D01 , cmd_R51_D08 , cmd_R53_D08 , cmd_R54_D08 , cmd_R64_D08 , cmd_R49_D08 , cmd_R35_D08 , cmd_R34_D05 , cmd_R35_D05 , cmd_R36_D05 , cmd_R51_D05 , cmd_R64_D05 , cmd_R65_D05 , cmd_R49_D05 , cmd_R4_D05 , cmd_R30_D05 , cmd_R4_D18 , cmd_R65_D18 , cmd_R66_D18 , cmd_R67_D18 , cmd_R36_D18 , cmd_R80_D18 , cmd_R79_Sw01 , cmd_R80_Sw01 , cmd_R81_Sw01 , cmd_R84_Sw01 , cmd_R66_Sw01 , cmd_R33_Sw01 , cmd_R55_D10 , cmd_R57_D10 , cmd_R58_D10 , cmd_R77_D10 , cmd_R69_D10 , cmd_R70_D10 , cmd_R6_D10 , cmd_R7_D10 , cmd_R38_D10 , cmd_R26_D09 , cmd_R37_D09 , cmd_R38_D09 , cmd_R55_D09 , cmd_R77_D09 , cmd_R69_D09 , cmd_R70_D09 , cmd_R6_D09 , cmd_R7_D09 , cmd_R8_D09 , cmd_R32_D09 , cmd_R28_D09 , cmd_R8_D20 , cmd_R28_D20 , cmd_R75_D20 , cmd_R76_D20 , cmd_R68_D20 , cmd_R37_D20 , cmd_R27_D23 , cmd_R68_D23 , cmd_R69_D23 , cmd_R70_D23 , cmd_R71_D23 , cmd_R73_D23 , cmd_R57_D23 , cmd_R76_D23 , cmd_R10_D23 , cmd_R16_D23 , cmd_R56_D23 , cmd_R41_D03 , cmd_R43_D03 , cmd_R44_D03 , cmd_R60_D03 , cmd_R39_D03 , cmd_R46_D03 , cmd_R2_D14 , cmd_R22_D14 , cmd_R61_D14 , cmd_R62_D14 , cmd_R40_D14 , cmd_R88_D14 , cmd_R21_Sw04 , cmd_R87_Sw04 , cmd_R88_Sw04 , cmd_R89_Sw04 , cmd_R61_Sw04 , cmd_R31_Sw04 , cmd_R11_D04 , cmd_R42_D04 , cmd_R45_D04 , cmd_R46_D04 , cmd_R47_D04 , cmd_R43_D04 , cmd_R44_D04 , cmd_R85_D04 , cmd_R89_D04 , cmd_R85_Sw03 , cmd_R86_Sw03 , cmd_R87_Sw03 , cmd_R89_Sw03 , cmd_R45_Sw03 , cmd_R31_Sw03 , cmd_R11_Sw03 , cmd_R42_Sw03 , cmd_R2_D15 , cmd_R3_D15 , cmd_R12_D15 , cmd_R62_D15 , cmd_R11_Sw02 , cmd_R42_Sw02 , cmd_R59_Sw02 , cmd_R60_Sw02 , cmd_R44_Sw02 , cmd_R47_Sw02 , cmd_R13_D07 , cmd_R48_D07 , cmd_R49_D07 , cmd_R50_D07 , cmd_R52_D07 , cmd_R53_D07 , cmd_R54_D07 , cmd_R81_D07 , cmd_R82_D07 , cmd_R81_Sw05 , cmd_R82_Sw05 , cmd_R83_Sw05 , cmd_R84_Sw05 , cmd_R48_Sw05 , cmd_R33_Sw05 , cmd_R13_Sw05 , cmd_R52_Sw05 , cmd_R13_D16 , cmd_R52_D16 , cmd_R63_D16 , cmd_R64_D16 , cmd_R54_D16 , cmd_R50_D16 , cmd_R4_D19 , cmd_R5_D19 , cmd_R14_D19 , cmd_R67_D19 , cmd_R8_D21 , cmd_R9_D21 , cmd_R15_D21 , cmd_R75_D21 , cmd_R37_D21 , cmd_R16_D24 , cmd_R56_D24 , cmd_R77_D24 , cmd_R78_D24 , cmd_R58_D24 , cmd_R69_D24 , cmd_R6_D24 : routeCommands := RELEASE;
	signal cmd_R6_D12 , cmd_R7_D12 , cmd_R69_D12 , cmd_R70_D12 , cmd_R71_D12 , cmd_R72_D12 , cmd_R73_D12 , cmd_R74_D12 : routeCommands := RELEASE;
	signal cmd_R1_T02 , cmd_R2_T04 , cmd_R3_T04 , cmd_R4_T06 , cmd_R5_T06 , cmd_R6_T08 , cmd_R7_T08 , cmd_R8_T10 , cmd_R9_T10 , cmd_R10_T12 , cmd_R11_T14 , cmd_R12_T16 , cmd_R13_T18 , cmd_R14_T20 , cmd_R15_T22 , cmd_R16_T24 , cmd_R17_L29 , cmd_R18_L30 , cmd_R19_L31 , cmd_R20_J35 , cmd_R21_J36 , cmd_R22_J37 , cmd_R23_J38 , cmd_R24_J40 , cmd_R25_J43 , cmd_R26_J45 , cmd_R27_J46 , cmd_R28_J47 , cmd_R29_J48 , cmd_R30_X50 , cmd_R31_X51 , cmd_R32_X52 , cmd_R33_X53 , cmd_R34_C54 , cmd_R35_S55 , cmd_R36_S55 , cmd_R37_S59 , cmd_R38_S59 , cmd_R39_S64 , cmd_R40_S64 , cmd_R41_C67 , cmd_R42_B68 , cmd_R43_S69 , cmd_R44_S69 , cmd_R45_C70 , cmd_R46_S71 , cmd_R47_S71 , cmd_R48_C73 , cmd_R49_S74 , cmd_R50_S74 , cmd_R51_C76 , cmd_R52_B77 , cmd_R53_S78 , cmd_R54_S78 , cmd_R55_C79 , cmd_R56_B80 , cmd_R57_S81 , cmd_R58_S81 , cmd_R59_S84 , cmd_R60_S84 , cmd_R61_S86 , cmd_R62_S86 , cmd_R63_S93 , cmd_R64_S93 , cmd_R65_C94 , cmd_R66_S95 , cmd_R67_S95 , cmd_R68_S101 , cmd_R69_S101 , cmd_R70_S101 , cmd_R71_S104 , cmd_R72_S104 , cmd_R73_S107 , cmd_R74_S107 , cmd_R75_S110 , cmd_R76_S110 , cmd_R77_S117 , cmd_R78_S117 , cmd_R79_C119 , cmd_R80_S120 , cmd_R81_S120 , cmd_R82_C122 , cmd_R83_S123 , cmd_R84_S123 , cmd_R85_C125 , cmd_R86_S126 , cmd_R87_S126 , cmd_R88_S129 , cmd_R89_S129 : routeCommands := RELEASE;
	signal cmd_R1_S64 , cmd_R2_J35 , cmd_R3_T15 , cmd_R4_C54 , cmd_R5_T19 , cmd_R6_S117 , cmd_R7_C79 , cmd_R8_J45 , cmd_R9_T21 , cmd_R10_S101 , cmd_R11_S126 , cmd_R12_T03 , cmd_R13_S123 , cmd_R14_T05 , cmd_R15_T09 , cmd_R16_S104 , cmd_R17_J48 , cmd_R18_X50 , cmd_R19_X52 , cmd_R20_T01 , cmd_R21_J38 , cmd_R22_J35 , cmd_R23_L30 , cmd_R24_L31 , cmd_R25_X53 , cmd_R26_J43 , cmd_R27_L29 , cmd_R28_J45 , cmd_R29_T11 , cmd_R30_S55 , cmd_R31_S129 , cmd_R32_S59 , cmd_R33_S120 , cmd_R34_X51 , cmd_R35_S78 , cmd_R36_S95 , cmd_R37_S110 , cmd_R38_S81 , cmd_R39_S69 , cmd_R40_S86 , cmd_R41_T01 , cmd_R42_S126 , cmd_R43_C70 , cmd_R44_B68 , cmd_R45_S126 , cmd_R46_C67 , cmd_R47_S84 , cmd_R48_S123 , cmd_R49_C76 , cmd_R50_S93 , cmd_R51_X51 , cmd_R52_S123 , cmd_R53_C73 , cmd_R54_B77 , cmd_R55_J43 , cmd_R56_S104 , cmd_R57_S107 , cmd_R58_B80 , cmd_R59_T13 , cmd_R60_T01 , cmd_R61_J36 , cmd_R62_T03 , cmd_R63_T17 , cmd_R64_X51 , cmd_R65_C54 , cmd_R66_C119 , cmd_R67_T05 , cmd_R68_J47 , cmd_R69_S117 , cmd_R70_C79 , cmd_R71_L29 , cmd_R72_T07 , cmd_R73_L29 , cmd_R74_T07 , cmd_R75_T09 , cmd_R76_J46 , cmd_R77_J43 , cmd_R78_T23 , cmd_R79_J40 , cmd_R80_C94 , cmd_R81_S74 , cmd_R82_S74 , cmd_R83_T25 , cmd_R84_J40 , cmd_R85_S71 , cmd_R86_T27 , cmd_R87_J38 , cmd_R88_J37 , cmd_R89_S71 : routeCommands := RELEASE;
begin
	levelCrossing_Lc01 : levelCrossing_0 port map(track_ne98 => tracks_i(20), track_ne996 => tracks_i(45), track_ne99 => tracks_i(21), R30_command => cmd_R30_Lc01, R31_command => cmd_R31_Lc01, R34_command => cmd_R34_Lc01, R51_command => cmd_R51_Lc01, R64_command => cmd_R64_Lc01, indication => levelCrossings_i(0), command  => levelCrossings_o(0), correspondence => state_Lc01, clock => clock, reset => reset);
	levelCrossing_Lc04 : levelCrossing_1 port map(track_ne100 => tracks_i(22), track_ne992 => tracks_i(41), track_ne101 => tracks_i(23), R32_command => cmd_R32_Lc04, R33_command => cmd_R33_Lc04, indication => levelCrossings_i(1), command  => levelCrossings_o(1), correspondence => state_Lc04, clock => clock, reset => reset);
	singleSwitch_D01 : singleSwitch_0 port map(R20_command => cmd_R20_D01, R39_command => cmd_R39_D01, R40_command => cmd_R40_D01, R41_command => cmd_R41_D01, R60_command => cmd_R60_D01, R1_command => cmd_R1_D01, R22_command => cmd_R22_D01, R46_command => cmd_R46_D01, R2_command => cmd_R2_D01, indication => singleSwitches_i(0), command => singleSwitches_o(0), correspondence => state_D01, clock => clock, reset => reset);
	singleSwitch_D08 : singleSwitch_1 port map(R51_command => cmd_R51_D08, R53_command => cmd_R53_D08, R54_command => cmd_R54_D08, R64_command => cmd_R64_D08, R49_command => cmd_R49_D08, R35_command => cmd_R35_D08, indication => singleSwitches_i(1), command => singleSwitches_o(1), correspondence => state_D08, clock => clock, reset => reset);
	singleSwitch_D05 : singleSwitch_2 port map(R34_command => cmd_R34_D05, R35_command => cmd_R35_D05, R36_command => cmd_R36_D05, R51_command => cmd_R51_D05, R64_command => cmd_R64_D05, R65_command => cmd_R65_D05, R49_command => cmd_R49_D05, R4_command => cmd_R4_D05, R30_command => cmd_R30_D05, indication => singleSwitches_i(2), command => singleSwitches_o(2), correspondence => state_D05, clock => clock, reset => reset);
	singleSwitch_D18 : singleSwitch_3 port map(R4_command => cmd_R4_D18, R65_command => cmd_R65_D18, R66_command => cmd_R66_D18, R67_command => cmd_R67_D18, R36_command => cmd_R36_D18, R80_command => cmd_R80_D18, indication => singleSwitches_i(3), command => singleSwitches_o(3), correspondence => state_D18, clock => clock, reset => reset);
	singleSwitch_Sw01 : singleSwitch_4 port map(R79_command => cmd_R79_Sw01, R80_command => cmd_R80_Sw01, R81_command => cmd_R81_Sw01, R84_command => cmd_R84_Sw01, R66_command => cmd_R66_Sw01, R33_command => cmd_R33_Sw01, indication => singleSwitches_i(4), command => singleSwitches_o(4), correspondence => state_Sw01, clock => clock, reset => reset);
	singleSwitch_D10 : singleSwitch_5 port map(R55_command => cmd_R55_D10, R57_command => cmd_R57_D10, R58_command => cmd_R58_D10, R77_command => cmd_R77_D10, R69_command => cmd_R69_D10, R70_command => cmd_R70_D10, R6_command => cmd_R6_D10, R7_command => cmd_R7_D10, R38_command => cmd_R38_D10, indication => singleSwitches_i(5), command => singleSwitches_o(5), correspondence => state_D10, clock => clock, reset => reset);
	singleSwitch_D09 : singleSwitch_6 port map(R26_command => cmd_R26_D09, R37_command => cmd_R37_D09, R38_command => cmd_R38_D09, R55_command => cmd_R55_D09, R77_command => cmd_R77_D09, R69_command => cmd_R69_D09, R70_command => cmd_R70_D09, R6_command => cmd_R6_D09, R7_command => cmd_R7_D09, R8_command => cmd_R8_D09, R32_command => cmd_R32_D09, R28_command => cmd_R28_D09, indication => singleSwitches_i(6), command => singleSwitches_o(6), correspondence => state_D09, clock => clock, reset => reset);
	singleSwitch_D20 : singleSwitch_7 port map(R8_command => cmd_R8_D20, R28_command => cmd_R28_D20, R75_command => cmd_R75_D20, R76_command => cmd_R76_D20, R68_command => cmd_R68_D20, R37_command => cmd_R37_D20, indication => singleSwitches_i(7), command => singleSwitches_o(7), correspondence => state_D20, clock => clock, reset => reset);
	singleSwitch_D23 : singleSwitch_8 port map(R27_command => cmd_R27_D23, R68_command => cmd_R68_D23, R69_command => cmd_R69_D23, R70_command => cmd_R70_D23, R71_command => cmd_R71_D23, R73_command => cmd_R73_D23, R57_command => cmd_R57_D23, R76_command => cmd_R76_D23, R10_command => cmd_R10_D23, R16_command => cmd_R16_D23, R56_command => cmd_R56_D23, indication => singleSwitches_i(8), command => singleSwitches_o(8), correspondence => state_D23, clock => clock, reset => reset);
	singleSwitch_D03 : singleSwitch_9 port map(R41_command => cmd_R41_D03, R43_command => cmd_R43_D03, R44_command => cmd_R44_D03, R60_command => cmd_R60_D03, R39_command => cmd_R39_D03, R46_command => cmd_R46_D03, indication => singleSwitches_i(9), command => singleSwitches_o(9), correspondence => state_D03, clock => clock, reset => reset);
	singleSwitch_D14 : singleSwitch_10 port map(R2_command => cmd_R2_D14, R22_command => cmd_R22_D14, R61_command => cmd_R61_D14, R62_command => cmd_R62_D14, R40_command => cmd_R40_D14, R88_command => cmd_R88_D14, indication => singleSwitches_i(10), command => singleSwitches_o(10), correspondence => state_D14, clock => clock, reset => reset);
	singleSwitch_Sw04 : singleSwitch_11 port map(R21_command => cmd_R21_Sw04, R87_command => cmd_R87_Sw04, R88_command => cmd_R88_Sw04, R89_command => cmd_R89_Sw04, R61_command => cmd_R61_Sw04, R31_command => cmd_R31_Sw04, indication => singleSwitches_i(11), command => singleSwitches_o(11), correspondence => state_Sw04, clock => clock, reset => reset);
	singleSwitch_D04 : singleSwitch_12 port map(R11_command => cmd_R11_D04, R42_command => cmd_R42_D04, R45_command => cmd_R45_D04, R46_command => cmd_R46_D04, R47_command => cmd_R47_D04, R43_command => cmd_R43_D04, R44_command => cmd_R44_D04, R85_command => cmd_R85_D04, R89_command => cmd_R89_D04, indication => singleSwitches_i(12), command => singleSwitches_o(12), correspondence => state_D04, clock => clock, reset => reset);
	singleSwitch_Sw03 : singleSwitch_13 port map(R85_command => cmd_R85_Sw03, R86_command => cmd_R86_Sw03, R87_command => cmd_R87_Sw03, R89_command => cmd_R89_Sw03, R45_command => cmd_R45_Sw03, R31_command => cmd_R31_Sw03, R11_command => cmd_R11_Sw03, R42_command => cmd_R42_Sw03, indication => singleSwitches_i(13), command => singleSwitches_o(13), correspondence => state_Sw03, clock => clock, reset => reset);
	singleSwitch_D15 : singleSwitch_14 port map(R2_command => cmd_R2_D15, R3_command => cmd_R3_D15, R12_command => cmd_R12_D15, R62_command => cmd_R62_D15, indication => singleSwitches_i(14), command => singleSwitches_o(14), correspondence => state_D15, clock => clock, reset => reset);
	singleSwitch_Sw02 : singleSwitch_15 port map(R11_command => cmd_R11_Sw02, R42_command => cmd_R42_Sw02, R59_command => cmd_R59_Sw02, R60_command => cmd_R60_Sw02, R44_command => cmd_R44_Sw02, R47_command => cmd_R47_Sw02, indication => singleSwitches_i(15), command => singleSwitches_o(15), correspondence => state_Sw02, clock => clock, reset => reset);
	singleSwitch_D07 : singleSwitch_16 port map(R13_command => cmd_R13_D07, R48_command => cmd_R48_D07, R49_command => cmd_R49_D07, R50_command => cmd_R50_D07, R52_command => cmd_R52_D07, R53_command => cmd_R53_D07, R54_command => cmd_R54_D07, R81_command => cmd_R81_D07, R82_command => cmd_R82_D07, indication => singleSwitches_i(16), command => singleSwitches_o(16), correspondence => state_D07, clock => clock, reset => reset);
	singleSwitch_Sw05 : singleSwitch_17 port map(R81_command => cmd_R81_Sw05, R82_command => cmd_R82_Sw05, R83_command => cmd_R83_Sw05, R84_command => cmd_R84_Sw05, R48_command => cmd_R48_Sw05, R33_command => cmd_R33_Sw05, R13_command => cmd_R13_Sw05, R52_command => cmd_R52_Sw05, indication => singleSwitches_i(17), command => singleSwitches_o(17), correspondence => state_Sw05, clock => clock, reset => reset);
	singleSwitch_D16 : singleSwitch_18 port map(R13_command => cmd_R13_D16, R52_command => cmd_R52_D16, R63_command => cmd_R63_D16, R64_command => cmd_R64_D16, R54_command => cmd_R54_D16, R50_command => cmd_R50_D16, indication => singleSwitches_i(18), command => singleSwitches_o(18), correspondence => state_D16, clock => clock, reset => reset);
	singleSwitch_D19 : singleSwitch_19 port map(R4_command => cmd_R4_D19, R5_command => cmd_R5_D19, R14_command => cmd_R14_D19, R67_command => cmd_R67_D19, indication => singleSwitches_i(19), command => singleSwitches_o(19), correspondence => state_D19, clock => clock, reset => reset);
	singleSwitch_D21 : singleSwitch_20 port map(R8_command => cmd_R8_D21, R9_command => cmd_R9_D21, R15_command => cmd_R15_D21, R75_command => cmd_R75_D21, R37_command => cmd_R37_D21, indication => singleSwitches_i(20), command => singleSwitches_o(20), correspondence => state_D21, clock => clock, reset => reset);
	singleSwitch_D24 : singleSwitch_21 port map(R16_command => cmd_R16_D24, R56_command => cmd_R56_D24, R77_command => cmd_R77_D24, R78_command => cmd_R78_D24, R58_command => cmd_R58_D24, R69_command => cmd_R69_D24, R6_command => cmd_R6_D24, indication => singleSwitches_i(21), command => singleSwitches_o(21), correspondence => state_D24, clock => clock, reset => reset);
	doubleSwitch_D12 : doubleSwitch_0 port map(R6_command => cmd_R6_D12, R7_command => cmd_R7_D12, R69_command => cmd_R69_D12, R70_command => cmd_R70_D12, R71_command => cmd_R71_D12, R72_command => cmd_R72_D12, R73_command => cmd_R73_D12, R74_command => cmd_R74_D12, indication => doubleSwitches_i, command => doubleSwitches_o, correspondence=> state_D12, clock => clock, reset => reset);
	railwaySignal_T01 : railwaySignal_0 port map(R20_command => cmd_R20_T01, R41_command => cmd_R41_T01, R60_command => cmd_R60_T01, track_ne991 => tracks_i(0), indication => signals_i(0), command => signals_o(0), correspondence_T01 => state_T01, clock => clock, reset => reset);
	railwaySignal_T02 : railwaySignal_1 port map(R1_command => cmd_R1_T02, track_ne991 => tracks_i(0), track_ne290 => tracks_i(8), track_ne288 => tracks_i(7), correspondence_S64 => state_S64, correspondence_S69 => state_S69, correspondence_S86 => state_S86, D01_state => state_D01, indication => signals_i(1), command => signals_o(1), correspondence_T02 => state_T02, clock => clock, reset => reset);
	railwaySignal_S64 : railwaySignal_2 port map(R39_command => cmd_R39_S64, R40_command => cmd_R40_S64, R1_command => cmd_R1_S64, track_ne991 => tracks_i(0), track_ne288 => tracks_i(7), track_ne290 => tracks_i(8), track_ne295 => tracks_i(10), track_ne110 => tracks_i(26), track_ne292 => tracks_i(9), track_ne111 => tracks_i(27), track_ne377 => tracks_i(12), correspondence_S69 => state_S69, correspondence_S86 => state_S86, correspondence_C70 => state_C70, correspondence_B68 => state_B68, correspondence_J36 => state_J36, correspondence_T03 => state_T03, D01_state => state_D01, D03_state => state_D03, D14_state => state_D14, D15_state => state_D15, indication => signals_i(2), command => signals_o(2), correspondence_S64 => state_S64, clock => clock, reset => reset);
	railwaySignal_S78 : railwaySignal_3 port map(R53_command => cmd_R53_S78, R54_command => cmd_R54_S78, R35_command => cmd_R35_S78, track_ne61 => tracks_i(1), track_ne404 => tracks_i(15), track_ne123 => tracks_i(30), track_ne400 => tracks_i(14), track_ne407 => tracks_i(16), correspondence_C73 => state_C73, correspondence_B77 => state_B77, correspondence_S123 => state_S123, D08_state => state_D08, D07_state => state_D07, D16_state => state_D16, indication => signals_i(3), command => signals_o(3), correspondence_S78 => state_S78, clock => clock, reset => reset);
	railwaySignal_C54 : railwaySignal_4 port map(R34_command => cmd_R34_C54, R4_command => cmd_R4_C54, R65_command => cmd_R65_C54, track_ne63 => tracks_i(2), track_ne99 => tracks_i(21), track_ne98 => tracks_i(20), track_ne996 => tracks_i(45), correspondence_X51 => state_X51, correspondence_S129 => state_S129, D05_state => state_D05, Lc01_state => state_Lc01, indication => signals_i(4), command => signals_o(4), correspondence_C54 => state_C54, clock => clock, reset => reset);
	railwaySignal_S95 : railwaySignal_5 port map(R66_command => cmd_R66_S95, R67_command => cmd_R67_S95, R36_command => cmd_R36_S95, track_ne63 => tracks_i(2), track_ne65 => tracks_i(3), track_ne124 => tracks_i(31), track_ne421 => tracks_i(17), track_ne992 => tracks_i(41), correspondence_C119 => state_C119, correspondence_T05 => state_T05, correspondence_J40 => state_J40, D18_state => state_D18, Sw01_state => state_Sw01, D19_state => state_D19, indication => signals_i(5), command => signals_o(5), correspondence_S95 => state_S95, clock => clock, reset => reset);
	railwaySignal_C94 : railwaySignal_6 port map(R65_command => cmd_R65_C94, R80_command => cmd_R80_C94, track_ne65 => tracks_i(3), track_ne63 => tracks_i(2), track_ne98 => tracks_i(20), track_ne99 => tracks_i(21), correspondence_C54 => state_C54, correspondence_X51 => state_X51, D18_state => state_D18, D05_state => state_D05, indication => signals_i(6), command => signals_o(6), correspondence_C94 => state_C94, clock => clock, reset => reset);
	railwaySignal_C119 : railwaySignal_7 port map(R79_command => cmd_R79_C119, R66_command => cmd_R66_C119, track_ne65 => tracks_i(3), track_ne992 => tracks_i(41), track_ne100 => tracks_i(22), correspondence_J40 => state_J40, correspondence_L31 => state_L31, Sw01_state => state_Sw01, indication => signals_i(7), command => signals_o(7), correspondence_C119 => state_C119, clock => clock, reset => reset);
	railwaySignal_S81 : railwaySignal_8 port map(R57_command => cmd_R57_S81, R58_command => cmd_R58_S81, R38_command => cmd_R38_S81, track_ne910 => tracks_i(4), track_ne130 => tracks_i(35), track_ne135 => tracks_i(40), track_ne129 => tracks_i(34), track_ne450 => tracks_i(18), track_ne114 => tracks_i(6), track_ne127 => tracks_i(33), correspondence_S107 => state_S107, correspondence_B80 => state_B80, correspondence_L29 => state_L29, correspondence_T07 => state_T07, correspondence_S104 => state_S104, D10_state => state_D10, D23_state => state_D23, D12_state => state_D12, D24_state => state_D24, indication => signals_i(8), command => signals_o(8), correspondence_S81 => state_S81, clock => clock, reset => reset);
	railwaySignal_J45 : railwaySignal_9 port map(R26_command => cmd_R26_J45, R8_command => cmd_R8_J45, R28_command => cmd_R28_J45, track_ne912 => tracks_i(5), track_ne101 => tracks_i(23), track_ne100 => tracks_i(22), correspondence_J43 => state_J43, correspondence_X53 => state_X53, D09_state => state_D09, indication => signals_i(9), command => signals_o(9), correspondence_J45 => state_J45, clock => clock, reset => reset);
	railwaySignal_S110 : railwaySignal_10 port map(R75_command => cmd_R75_S110, R76_command => cmd_R76_S110, R37_command => cmd_R37_S110, track_ne912 => tracks_i(5), track_ne131 => tracks_i(36), track_ne465 => tracks_i(19), track_ne132 => tracks_i(37), track_ne114 => tracks_i(6), correspondence_T09 => state_T09, correspondence_J46 => state_J46, correspondence_L29 => state_L29, D20_state => state_D20, D21_state => state_D21, D23_state => state_D23, indication => signals_i(10), command => signals_o(10), correspondence_S110 => state_S110, clock => clock, reset => reset);
	railwaySignal_L29 : railwaySignal_11 port map(R17_command => cmd_R17_L29, R27_command => cmd_R27_L29, R71_command => cmd_R71_L29, R73_command => cmd_R73_L29, track_ne114 => tracks_i(6), track_ne102 => tracks_i(24), correspondence_J48 => state_J48, correspondence_T11 => state_T11, indication => signals_i(11), command => signals_o(11), correspondence_L29 => state_L29, clock => clock, reset => reset);
	railwaySignal_J48 : railwaySignal_12 port map(R29_command => cmd_R29_J48, R17_command => cmd_R17_J48, track_ne114 => tracks_i(6), track_ne102 => tracks_i(24), correspondence_T11 => state_T11, indication => signals_i(12), command => signals_o(12), correspondence_J48 => state_J48, clock => clock, reset => reset);
	railwaySignal_S101 : railwaySignal_13 port map(R68_command => cmd_R68_S101, R69_command => cmd_R69_S101, R70_command => cmd_R70_S101, R10_command => cmd_R10_S101, track_ne114 => tracks_i(6), track_ne132 => tracks_i(37), track_ne129 => tracks_i(34), track_ne127 => tracks_i(33), track_ne130 => tracks_i(35), track_ne912 => tracks_i(5), track_ne910 => tracks_i(4), track_ne134 => tracks_i(39), track_ne135 => tracks_i(40), track_ne101 => tracks_i(23), correspondence_J47 => state_J47, correspondence_S117 => state_S117, correspondence_C79 => state_C79, correspondence_J45 => state_J45, correspondence_J43 => state_J43, correspondence_T23 => state_T23, D23_state => state_D23, D20_state => state_D20, D12_state => state_D12, D09_state => state_D09, D10_state => state_D10, D24_state => state_D24, indication => signals_i(13), command => signals_o(13), correspondence_S101 => state_S101, clock => clock, reset => reset);
	railwaySignal_S69 : railwaySignal_14 port map(R43_command => cmd_R43_S69, R44_command => cmd_R44_S69, R39_command => cmd_R39_S69, track_ne288 => tracks_i(7), track_ne295 => tracks_i(10), track_ne110 => tracks_i(26), track_ne297 => tracks_i(11), track_ne384 => tracks_i(13), correspondence_C70 => state_C70, correspondence_B68 => state_B68, correspondence_S126 => state_S126, D03_state => state_D03, D04_state => state_D04, Sw02_state => state_Sw02, indication => signals_i(14), command => signals_o(14), correspondence_S69 => state_S69, clock => clock, reset => reset);
	railwaySignal_J35 : railwaySignal_15 port map(R20_command => cmd_R20_J35, R2_command => cmd_R2_J35, R22_command => cmd_R22_J35, track_ne290 => tracks_i(8), track_ne991 => tracks_i(0), correspondence_T01 => state_T01, D01_state => state_D01, indication => signals_i(15), command => signals_o(15), correspondence_J35 => state_J35, clock => clock, reset => reset);
	railwaySignal_S86 : railwaySignal_16 port map(R61_command => cmd_R61_S86, R62_command => cmd_R62_S86, R40_command => cmd_R40_S86, track_ne290 => tracks_i(8), track_ne292 => tracks_i(9), track_ne111 => tracks_i(27), track_ne377 => tracks_i(12), track_ne996 => tracks_i(45), correspondence_J36 => state_J36, correspondence_T03 => state_T03, correspondence_J38 => state_J38, D14_state => state_D14, Sw04_state => state_Sw04, D15_state => state_D15, indication => signals_i(16), command => signals_o(16), correspondence_S86 => state_S86, clock => clock, reset => reset);
	railwaySignal_J36 : railwaySignal_17 port map(R21_command => cmd_R21_J36, R61_command => cmd_R61_J36, track_ne292 => tracks_i(9), track_ne996 => tracks_i(45), track_ne98 => tracks_i(20), correspondence_J38 => state_J38, correspondence_L30 => state_L30, Sw04_state => state_Sw04, indication => signals_i(17), command => signals_o(17), correspondence_J36 => state_J36, clock => clock, reset => reset);
	railwaySignal_J37 : railwaySignal_18 port map(R22_command => cmd_R22_J37, R88_command => cmd_R88_J37, track_ne292 => tracks_i(9), track_ne290 => tracks_i(8), track_ne991 => tracks_i(0), correspondence_J35 => state_J35, correspondence_T01 => state_T01, D14_state => state_D14, D01_state => state_D01, indication => signals_i(18), command => signals_o(18), correspondence_J37 => state_J37, clock => clock, reset => reset);
	railwaySignal_C67 : railwaySignal_19 port map(R41_command => cmd_R41_C67, R46_command => cmd_R46_C67, track_ne295 => tracks_i(10), track_ne288 => tracks_i(7), track_ne991 => tracks_i(0), correspondence_T01 => state_T01, D01_state => state_D01, D03_state => state_D03, indication => signals_i(19), command => signals_o(19), correspondence_C67 => state_C67, clock => clock, reset => reset);
	railwaySignal_C70 : railwaySignal_20 port map(R45_command => cmd_R45_C70, R43_command => cmd_R43_C70, track_ne295 => tracks_i(10), track_ne297 => tracks_i(11), track_ne996 => tracks_i(45), track_ne997 => tracks_i(46), track_ne995 => tracks_i(44), correspondence_S126 => state_S126, correspondence_T27 => state_T27, correspondence_J38 => state_J38, D04_state => state_D04, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication => signals_i(20), command => signals_o(20), correspondence_C70 => state_C70, clock => clock, reset => reset);
	railwaySignal_S71 : railwaySignal_21 port map(R46_command => cmd_R46_S71, R47_command => cmd_R47_S71, R85_command => cmd_R85_S71, R89_command => cmd_R89_S71, track_ne297 => tracks_i(11), track_ne295 => tracks_i(10), track_ne384 => tracks_i(13), track_ne991 => tracks_i(0), track_ne288 => tracks_i(7), track_ne104 => tracks_i(25), track_ne110 => tracks_i(26), correspondence_C67 => state_C67, correspondence_S84 => state_S84, correspondence_T01 => state_T01, correspondence_T13 => state_T13, D04_state => state_D04, D01_state => state_D01, D03_state => state_D03, Sw02_state => state_Sw02, indication => signals_i(21), command => signals_o(21), correspondence_S71 => state_S71, clock => clock, reset => reset);
	railwaySignal_S126 : railwaySignal_22 port map(R86_command => cmd_R86_S126, R87_command => cmd_R87_S126, R11_command => cmd_R11_S126, R42_command => cmd_R42_S126, R45_command => cmd_R45_S126, track_ne297 => tracks_i(11), track_ne995 => tracks_i(44), track_ne997 => tracks_i(46), track_ne996 => tracks_i(45), track_ne98 => tracks_i(20), correspondence_T27 => state_T27, correspondence_J38 => state_J38, correspondence_L30 => state_L30, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication => signals_i(22), command => signals_o(22), correspondence_S126 => state_S126, clock => clock, reset => reset);
	railwaySignal_T03 : railwaySignal_23 port map(R12_command => cmd_R12_T03, R62_command => cmd_R62_T03, track_ne377 => tracks_i(12), indication => signals_i(23), command => signals_o(23), correspondence_T03 => state_T03, clock => clock, reset => reset);
	railwaySignal_T04 : railwaySignal_24 port map(R2_command => cmd_R2_T04, R3_command => cmd_R3_T04, track_ne377 => tracks_i(12), track_ne111 => tracks_i(27), track_ne290 => tracks_i(8), track_ne113 => tracks_i(28), track_ne991 => tracks_i(0), correspondence_J35 => state_J35, correspondence_T15 => state_T15, correspondence_T01 => state_T01, D14_state => state_D14, D15_state => state_D15, D01_state => state_D01, indication => signals_i(24), command => signals_o(24), correspondence_T04 => state_T04, clock => clock, reset => reset);
	railwaySignal_S84 : railwaySignal_25 port map(R59_command => cmd_R59_S84, R60_command => cmd_R60_S84, R47_command => cmd_R47_S84, track_ne384 => tracks_i(13), track_ne104 => tracks_i(25), track_ne110 => tracks_i(26), track_ne288 => tracks_i(7), track_ne991 => tracks_i(0), correspondence_T13 => state_T13, correspondence_T01 => state_T01, Sw02_state => state_Sw02, D01_state => state_D01, D03_state => state_D03, indication => signals_i(25), command => signals_o(25), correspondence_S84 => state_S84, clock => clock, reset => reset);
	railwaySignal_S74 : railwaySignal_26 port map(R49_command => cmd_R49_S74, R50_command => cmd_R50_S74, R81_command => cmd_R81_S74, R82_command => cmd_R82_S74, track_ne400 => tracks_i(14), track_ne404 => tracks_i(15), track_ne407 => tracks_i(16), track_ne61 => tracks_i(1), track_ne98 => tracks_i(20), track_ne99 => tracks_i(21), track_ne122 => tracks_i(29), track_ne123 => tracks_i(30), correspondence_C76 => state_C76, correspondence_S93 => state_S93, correspondence_X51 => state_X51, correspondence_T17 => state_T17, D07_state => state_D07, D05_state => state_D05, D08_state => state_D08, D16_state => state_D16, indication => signals_i(26), command => signals_o(26), correspondence_S74 => state_S74, clock => clock, reset => reset);
	railwaySignal_S123 : railwaySignal_27 port map(R83_command => cmd_R83_S123, R84_command => cmd_R84_S123, R13_command => cmd_R13_S123, R48_command => cmd_R48_S123, R52_command => cmd_R52_S123, track_ne400 => tracks_i(14), track_ne993 => tracks_i(42), track_ne994 => tracks_i(43), track_ne992 => tracks_i(41), track_ne100 => tracks_i(22), correspondence_T25 => state_T25, correspondence_J40 => state_J40, correspondence_L31 => state_L31, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication => signals_i(27), command => signals_o(27), correspondence_S123 => state_S123, clock => clock, reset => reset);
	railwaySignal_C73 : railwaySignal_28 port map(R48_command => cmd_R48_C73, R53_command => cmd_R53_C73, track_ne404 => tracks_i(15), track_ne400 => tracks_i(14), track_ne994 => tracks_i(43), track_ne992 => tracks_i(41), track_ne993 => tracks_i(42), correspondence_S123 => state_S123, correspondence_T25 => state_T25, correspondence_J40 => state_J40, D07_state => state_D07, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication => signals_i(28), command => signals_o(28), correspondence_C73 => state_C73, clock => clock, reset => reset);
	railwaySignal_C76 : railwaySignal_29 port map(R51_command => cmd_R51_C76, R49_command => cmd_R49_C76, track_ne404 => tracks_i(15), track_ne61 => tracks_i(1), track_ne99 => tracks_i(21), track_ne98 => tracks_i(20), track_ne996 => tracks_i(45), correspondence_X51 => state_X51, correspondence_S129 => state_S129, D05_state => state_D05, D08_state => state_D08, Lc01_state => state_Lc01, indication => signals_i(29), command => signals_o(29), correspondence_C76 => state_C76, clock => clock, reset => reset);
	railwaySignal_S93 : railwaySignal_30 port map(R63_command => cmd_R63_S93, R64_command => cmd_R64_S93, R50_command => cmd_R50_S93, track_ne407 => tracks_i(16), track_ne122 => tracks_i(29), track_ne123 => tracks_i(30), track_ne61 => tracks_i(1), track_ne99 => tracks_i(21), track_ne98 => tracks_i(20), track_ne996 => tracks_i(45), correspondence_T17 => state_T17, correspondence_X51 => state_X51, correspondence_S129 => state_S129, D16_state => state_D16, D05_state => state_D05, D08_state => state_D08, Lc01_state => state_Lc01, indication => signals_i(30), command => signals_o(30), correspondence_S93 => state_S93, clock => clock, reset => reset);
	railwaySignal_T05 : railwaySignal_31 port map(R14_command => cmd_R14_T05, R67_command => cmd_R67_T05, track_ne421 => tracks_i(17), indication => signals_i(31), command => signals_o(31), correspondence_T05 => state_T05, clock => clock, reset => reset);
	railwaySignal_T06 : railwaySignal_32 port map(R4_command => cmd_R4_T06, R5_command => cmd_R5_T06, track_ne421 => tracks_i(17), track_ne124 => tracks_i(31), track_ne63 => tracks_i(2), track_ne126 => tracks_i(32), track_ne98 => tracks_i(20), track_ne99 => tracks_i(21), correspondence_C54 => state_C54, correspondence_T19 => state_T19, correspondence_X51 => state_X51, D18_state => state_D18, D19_state => state_D19, D05_state => state_D05, indication => signals_i(32), command => signals_o(32), correspondence_T06 => state_T06, clock => clock, reset => reset);
	railwaySignal_T07 : railwaySignal_33 port map(R72_command => cmd_R72_T07, R74_command => cmd_R74_T07, track_ne450 => tracks_i(18), indication => signals_i(33), command => signals_o(33), correspondence_T07 => state_T07, clock => clock, reset => reset);
	railwaySignal_T08 : railwaySignal_34 port map(R6_command => cmd_R6_T08, R7_command => cmd_R7_T08, track_ne450 => tracks_i(18), track_ne127 => tracks_i(33), track_ne130 => tracks_i(35), track_ne910 => tracks_i(4), track_ne134 => tracks_i(39), track_ne135 => tracks_i(40), track_ne101 => tracks_i(23), correspondence_S117 => state_S117, correspondence_C79 => state_C79, correspondence_J43 => state_J43, correspondence_T23 => state_T23, D12_state => state_D12, D09_state => state_D09, D10_state => state_D10, D24_state => state_D24, indication => signals_i(34), command => signals_o(34), correspondence_T08 => state_T08, clock => clock, reset => reset);
	railwaySignal_T09 : railwaySignal_35 port map(R15_command => cmd_R15_T09, R75_command => cmd_R75_T09, track_ne465 => tracks_i(19), indication => signals_i(35), command => signals_o(35), correspondence_T09 => state_T09, clock => clock, reset => reset);
	railwaySignal_T10 : railwaySignal_36 port map(R8_command => cmd_R8_T10, R9_command => cmd_R9_T10, track_ne465 => tracks_i(19), track_ne131 => tracks_i(36), track_ne912 => tracks_i(5), track_ne133 => tracks_i(38), track_ne101 => tracks_i(23), correspondence_J45 => state_J45, correspondence_T21 => state_T21, correspondence_J43 => state_J43, D20_state => state_D20, D21_state => state_D21, D09_state => state_D09, indication => signals_i(36), command => signals_o(36), correspondence_T10 => state_T10, clock => clock, reset => reset);
	railwaySignal_L30 : railwaySignal_37 port map(R18_command => cmd_R18_L30, R23_command => cmd_R23_L30, track_ne98 => tracks_i(20), track_ne99 => tracks_i(21), correspondence_X50 => state_X50, correspondence_S55 => state_S55, indication => signals_i(37), command => signals_o(37), correspondence_L30 => state_L30, clock => clock, reset => reset);
	railwaySignal_X50 : railwaySignal_38 port map(R30_command => cmd_R30_X50, R18_command => cmd_R18_X50, track_ne98 => tracks_i(20), track_ne99 => tracks_i(21), track_ne63 => tracks_i(2), track_ne61 => tracks_i(1), correspondence_S55 => state_S55, correspondence_S78 => state_S78, correspondence_S95 => state_S95, D05_state => state_D05, Lc01_state => state_Lc01, indication => signals_i(38), command => signals_o(38), correspondence_X50 => state_X50, clock => clock, reset => reset);
	railwaySignal_X51 : railwaySignal_39 port map(R31_command => cmd_R31_X51, R34_command => cmd_R34_X51, R51_command => cmd_R51_X51, R64_command => cmd_R64_X51, track_ne98 => tracks_i(20), track_ne996 => tracks_i(45), track_ne292 => tracks_i(9), track_ne997 => tracks_i(46), track_ne297 => tracks_i(11), correspondence_S129 => state_S129, correspondence_J37 => state_J37, correspondence_S71 => state_S71, Sw04_state => state_Sw04, Sw03_state => state_Sw03, Lc01_state => state_Lc01, indication => signals_i(39), command => signals_o(39), correspondence_X51 => state_X51, clock => clock, reset => reset);
	railwaySignal_S55 : railwaySignal_40 port map(R35_command => cmd_R35_S55, R36_command => cmd_R36_S55, R30_command => cmd_R30_S55, track_ne99 => tracks_i(21), track_ne61 => tracks_i(1), track_ne63 => tracks_i(2), track_ne404 => tracks_i(15), track_ne123 => tracks_i(30), track_ne421 => tracks_i(17), track_ne65 => tracks_i(3), track_ne124 => tracks_i(31), correspondence_S78 => state_S78, correspondence_S95 => state_S95, correspondence_C73 => state_C73, correspondence_B77 => state_B77, correspondence_C119 => state_C119, correspondence_T05 => state_T05, D05_state => state_D05, D08_state => state_D08, D18_state => state_D18, D19_state => state_D19, indication => signals_i(40), command => signals_o(40), correspondence_S55 => state_S55, clock => clock, reset => reset);
	railwaySignal_L31 : railwaySignal_41 port map(R19_command => cmd_R19_L31, R24_command => cmd_R24_L31, track_ne100 => tracks_i(22), track_ne101 => tracks_i(23), correspondence_X52 => state_X52, correspondence_S59 => state_S59, indication => signals_i(41), command => signals_o(41), correspondence_L31 => state_L31, clock => clock, reset => reset);
	railwaySignal_X52 : railwaySignal_42 port map(R32_command => cmd_R32_X52, R19_command => cmd_R19_X52, track_ne100 => tracks_i(22), track_ne101 => tracks_i(23), track_ne910 => tracks_i(4), track_ne912 => tracks_i(5), correspondence_S59 => state_S59, correspondence_S110 => state_S110, correspondence_S81 => state_S81, D09_state => state_D09, Lc04_state => state_Lc04, indication => signals_i(42), command => signals_o(42), correspondence_X52 => state_X52, clock => clock, reset => reset);
	railwaySignal_X53 : railwaySignal_43 port map(R33_command => cmd_R33_X53, R25_command => cmd_R25_X53, track_ne100 => tracks_i(22), track_ne992 => tracks_i(41), track_ne994 => tracks_i(43), track_ne65 => tracks_i(3), track_ne400 => tracks_i(14), correspondence_S120 => state_S120, correspondence_C94 => state_C94, correspondence_S74 => state_S74, Sw01_state => state_Sw01, Sw05_state => state_Sw05, Lc04_state => state_Lc04, indication => signals_i(43), command => signals_o(43), correspondence_X53 => state_X53, clock => clock, reset => reset);
	railwaySignal_J43 : railwaySignal_44 port map(R25_command => cmd_R25_J43, R26_command => cmd_R26_J43, R55_command => cmd_R55_J43, R77_command => cmd_R77_J43, track_ne101 => tracks_i(23), track_ne100 => tracks_i(22), track_ne992 => tracks_i(41), correspondence_X53 => state_X53, correspondence_S120 => state_S120, indication => signals_i(44), command => signals_o(44), correspondence_J43 => state_J43, clock => clock, reset => reset);
	railwaySignal_S59 : railwaySignal_45 port map(R37_command => cmd_R37_S59, R38_command => cmd_R38_S59, R32_command => cmd_R32_S59, track_ne101 => tracks_i(23), track_ne912 => tracks_i(5), track_ne910 => tracks_i(4), track_ne131 => tracks_i(36), track_ne132 => tracks_i(37), track_ne465 => tracks_i(19), track_ne130 => tracks_i(35), track_ne135 => tracks_i(40), correspondence_S110 => state_S110, correspondence_S81 => state_S81, correspondence_T09 => state_T09, correspondence_J46 => state_J46, correspondence_S107 => state_S107, correspondence_B80 => state_B80, D09_state => state_D09, D20_state => state_D20, D21_state => state_D21, D10_state => state_D10, indication => signals_i(45), command => signals_o(45), correspondence_S59 => state_S59, clock => clock, reset => reset);
	railwaySignal_T11 : railwaySignal_46 port map(R29_command => cmd_R29_T11, track_ne102 => tracks_i(24), indication => signals_i(46), command => signals_o(46), correspondence_T11 => state_T11, clock => clock, reset => reset);
	railwaySignal_T12 : railwaySignal_47 port map(R10_command => cmd_R10_T12, track_ne102 => tracks_i(24), track_ne114 => tracks_i(6), track_ne130 => tracks_i(35), track_ne129 => tracks_i(34), track_ne132 => tracks_i(37), track_ne127 => tracks_i(33), correspondence_S101 => state_S101, correspondence_J47 => state_J47, correspondence_S117 => state_S117, correspondence_C79 => state_C79, D23_state => state_D23, D12_state => state_D12, indication => signals_i(47), command => signals_o(47), correspondence_T12 => state_T12, clock => clock, reset => reset);
	railwaySignal_T13 : railwaySignal_48 port map(R59_command => cmd_R59_T13, track_ne104 => tracks_i(25), indication => signals_i(48), command => signals_o(48), correspondence_T13 => state_T13, clock => clock, reset => reset);
	railwaySignal_T14 : railwaySignal_49 port map(R11_command => cmd_R11_T14, track_ne104 => tracks_i(25), track_ne384 => tracks_i(13), track_ne297 => tracks_i(11), track_ne996 => tracks_i(45), track_ne997 => tracks_i(46), track_ne995 => tracks_i(44), correspondence_S126 => state_S126, correspondence_T27 => state_T27, correspondence_J38 => state_J38, D04_state => state_D04, Sw02_state => state_Sw02, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication => signals_i(49), command => signals_o(49), correspondence_T14 => state_T14, clock => clock, reset => reset);
	railwaySignal_B68 : railwaySignal_50 port map(R42_command => cmd_R42_B68, R44_command => cmd_R44_B68, track_ne110 => tracks_i(26), track_ne384 => tracks_i(13), track_ne297 => tracks_i(11), track_ne996 => tracks_i(45), track_ne997 => tracks_i(46), track_ne995 => tracks_i(44), correspondence_S126 => state_S126, correspondence_T27 => state_T27, correspondence_J38 => state_J38, D04_state => state_D04, Sw02_state => state_Sw02, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication => signals_i(50), command => signals_o(50), correspondence_B68 => state_B68, clock => clock, reset => reset);
	railwaySignal_T15 : railwaySignal_51 port map(R3_command => cmd_R3_T15, track_ne113 => tracks_i(28), indication => signals_i(51), command => signals_o(51), correspondence_T15 => state_T15, clock => clock, reset => reset);
	railwaySignal_T16 : railwaySignal_52 port map(R12_command => cmd_R12_T16, track_ne113 => tracks_i(28), track_ne377 => tracks_i(12), correspondence_T03 => state_T03, D15_state => state_D15, indication => signals_i(52), command => signals_o(52), correspondence_T16 => state_T16, clock => clock, reset => reset);
	railwaySignal_T17 : railwaySignal_53 port map(R63_command => cmd_R63_T17, track_ne122 => tracks_i(29), indication => signals_i(53), command => signals_o(53), correspondence_T17 => state_T17, clock => clock, reset => reset);
	railwaySignal_T18 : railwaySignal_54 port map(R13_command => cmd_R13_T18, track_ne122 => tracks_i(29), track_ne407 => tracks_i(16), track_ne400 => tracks_i(14), track_ne994 => tracks_i(43), track_ne992 => tracks_i(41), track_ne993 => tracks_i(42), correspondence_S123 => state_S123, correspondence_T25 => state_T25, correspondence_J40 => state_J40, D07_state => state_D07, D16_state => state_D16, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication => signals_i(54), command => signals_o(54), correspondence_T18 => state_T18, clock => clock, reset => reset);
	railwaySignal_B77 : railwaySignal_55 port map(R52_command => cmd_R52_B77, R54_command => cmd_R54_B77, track_ne123 => tracks_i(30), track_ne407 => tracks_i(16), track_ne400 => tracks_i(14), track_ne994 => tracks_i(43), track_ne992 => tracks_i(41), track_ne993 => tracks_i(42), correspondence_S123 => state_S123, correspondence_T25 => state_T25, correspondence_J40 => state_J40, D07_state => state_D07, D16_state => state_D16, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication => signals_i(55), command => signals_o(55), correspondence_B77 => state_B77, clock => clock, reset => reset);
	railwaySignal_T19 : railwaySignal_56 port map(R5_command => cmd_R5_T19, track_ne126 => tracks_i(32), indication => signals_i(56), command => signals_o(56), correspondence_T19 => state_T19, clock => clock, reset => reset);
	railwaySignal_T20 : railwaySignal_57 port map(R14_command => cmd_R14_T20, track_ne126 => tracks_i(32), track_ne421 => tracks_i(17), correspondence_T05 => state_T05, D19_state => state_D19, indication => signals_i(57), command => signals_o(57), correspondence_T20 => state_T20, clock => clock, reset => reset);
	railwaySignal_S104 : railwaySignal_58 port map(R71_command => cmd_R71_S104, R72_command => cmd_R72_S104, R16_command => cmd_R16_S104, R56_command => cmd_R56_S104, track_ne127 => tracks_i(33), track_ne129 => tracks_i(34), track_ne114 => tracks_i(6), track_ne450 => tracks_i(18), correspondence_L29 => state_L29, correspondence_T07 => state_T07, correspondence_J48 => state_J48, D23_state => state_D23, D12_state => state_D12, indication => signals_i(58), command => signals_o(58), correspondence_S104 => state_S104, clock => clock, reset => reset);
	railwaySignal_S117 : railwaySignal_59 port map(R77_command => cmd_R77_S117, R78_command => cmd_R78_S117, R6_command => cmd_R6_S117, R69_command => cmd_R69_S117, track_ne127 => tracks_i(33), track_ne135 => tracks_i(40), track_ne910 => tracks_i(4), track_ne101 => tracks_i(23), track_ne134 => tracks_i(39), track_ne100 => tracks_i(22), correspondence_J43 => state_J43, correspondence_T23 => state_T23, correspondence_X53 => state_X53, D09_state => state_D09, D10_state => state_D10, D24_state => state_D24, indication => signals_i(59), command => signals_o(59), correspondence_S117 => state_S117, clock => clock, reset => reset);
	railwaySignal_C79 : railwaySignal_60 port map(R55_command => cmd_R55_C79, R7_command => cmd_R7_C79, R70_command => cmd_R70_C79, track_ne130 => tracks_i(35), track_ne910 => tracks_i(4), track_ne101 => tracks_i(23), track_ne100 => tracks_i(22), correspondence_J43 => state_J43, correspondence_X53 => state_X53, D09_state => state_D09, D10_state => state_D10, indication => signals_i(60), command => signals_o(60), correspondence_C79 => state_C79, clock => clock, reset => reset);
	railwaySignal_S107 : railwaySignal_61 port map(R73_command => cmd_R73_S107, R74_command => cmd_R74_S107, R57_command => cmd_R57_S107, track_ne130 => tracks_i(35), track_ne129 => tracks_i(34), track_ne114 => tracks_i(6), track_ne450 => tracks_i(18), correspondence_L29 => state_L29, correspondence_T07 => state_T07, correspondence_J48 => state_J48, D23_state => state_D23, D12_state => state_D12, indication => signals_i(61), command => signals_o(61), correspondence_S107 => state_S107, clock => clock, reset => reset);
	railwaySignal_J46 : railwaySignal_62 port map(R27_command => cmd_R27_J46, R76_command => cmd_R76_J46, track_ne132 => tracks_i(37), track_ne114 => tracks_i(6), correspondence_L29 => state_L29, correspondence_J48 => state_J48, D23_state => state_D23, indication => signals_i(62), command => signals_o(62), correspondence_J46 => state_J46, clock => clock, reset => reset);
	railwaySignal_J47 : railwaySignal_63 port map(R28_command => cmd_R28_J47, R68_command => cmd_R68_J47, track_ne132 => tracks_i(37), track_ne912 => tracks_i(5), track_ne101 => tracks_i(23), correspondence_J45 => state_J45, correspondence_J43 => state_J43, D20_state => state_D20, D09_state => state_D09, indication => signals_i(63), command => signals_o(63), correspondence_J47 => state_J47, clock => clock, reset => reset);
	railwaySignal_T21 : railwaySignal_64 port map(R9_command => cmd_R9_T21, track_ne133 => tracks_i(38), indication => signals_i(64), command => signals_o(64), correspondence_T21 => state_T21, clock => clock, reset => reset);
	railwaySignal_T22 : railwaySignal_65 port map(R15_command => cmd_R15_T22, track_ne133 => tracks_i(38), track_ne465 => tracks_i(19), correspondence_T09 => state_T09, D21_state => state_D21, indication => signals_i(65), command => signals_o(65), correspondence_T22 => state_T22, clock => clock, reset => reset);
	railwaySignal_T23 : railwaySignal_66 port map(R78_command => cmd_R78_T23, track_ne134 => tracks_i(39), indication => signals_i(66), command => signals_o(66), correspondence_T23 => state_T23, clock => clock, reset => reset);
	railwaySignal_T24 : railwaySignal_67 port map(R16_command => cmd_R16_T24, track_ne134 => tracks_i(39), track_ne127 => tracks_i(33), track_ne129 => tracks_i(34), track_ne450 => tracks_i(18), track_ne114 => tracks_i(6), correspondence_S104 => state_S104, correspondence_L29 => state_L29, correspondence_T07 => state_T07, D24_state => state_D24, D23_state => state_D23, D12_state => state_D12, indication => signals_i(67), command => signals_o(67), correspondence_T24 => state_T24, clock => clock, reset => reset);
	railwaySignal_B80 : railwaySignal_68 port map(R56_command => cmd_R56_B80, R58_command => cmd_R58_B80, track_ne135 => tracks_i(40), track_ne127 => tracks_i(33), track_ne129 => tracks_i(34), track_ne450 => tracks_i(18), track_ne114 => tracks_i(6), correspondence_S104 => state_S104, correspondence_L29 => state_L29, correspondence_T07 => state_T07, D24_state => state_D24, D23_state => state_D23, D12_state => state_D12, indication => signals_i(68), command => signals_o(68), correspondence_B80 => state_B80, clock => clock, reset => reset);
	railwaySignal_J40 : railwaySignal_69 port map(R24_command => cmd_R24_J40, R79_command => cmd_R79_J40, R84_command => cmd_R84_J40, track_ne992 => tracks_i(41), track_ne100 => tracks_i(22), correspondence_L31 => state_L31, correspondence_X52 => state_X52, indication => signals_i(69), command => signals_o(69), correspondence_J40 => state_J40, clock => clock, reset => reset);
	railwaySignal_S120 : railwaySignal_70 port map(R80_command => cmd_R80_S120, R81_command => cmd_R81_S120, R33_command => cmd_R33_S120, track_ne992 => tracks_i(41), track_ne65 => tracks_i(3), track_ne994 => tracks_i(43), track_ne400 => tracks_i(14), track_ne63 => tracks_i(2), track_ne407 => tracks_i(16), track_ne404 => tracks_i(15), correspondence_C94 => state_C94, correspondence_S74 => state_S74, correspondence_C54 => state_C54, correspondence_C76 => state_C76, correspondence_S93 => state_S93, Sw01_state => state_Sw01, D18_state => state_D18, Sw05_state => state_Sw05, D07_state => state_D07, indication => signals_i(70), command => signals_o(70), correspondence_S120 => state_S120, clock => clock, reset => reset);
	railwaySignal_T25 : railwaySignal_71 port map(R83_command => cmd_R83_T25, track_ne993 => tracks_i(42), indication => signals_i(71), command => signals_o(71), correspondence_T25 => state_T25, clock => clock, reset => reset);
	railwaySignal_C122 : railwaySignal_72 port map(R82_command => cmd_R82_C122, track_ne993 => tracks_i(42), track_ne400 => tracks_i(14), track_ne407 => tracks_i(16), track_ne404 => tracks_i(15), correspondence_S74 => state_S74, correspondence_C76 => state_C76, correspondence_S93 => state_S93, Sw05_state => state_Sw05, D07_state => state_D07, indication => signals_i(72), command => signals_o(72), correspondence_C122 => state_C122, clock => clock, reset => reset);
	railwaySignal_T27 : railwaySignal_73 port map(R86_command => cmd_R86_T27, track_ne995 => tracks_i(44), indication => signals_i(73), command => signals_o(73), correspondence_T27 => state_T27, clock => clock, reset => reset);
	railwaySignal_C125 : railwaySignal_74 port map(R85_command => cmd_R85_C125, track_ne995 => tracks_i(44), track_ne297 => tracks_i(11), track_ne384 => tracks_i(13), track_ne295 => tracks_i(10), correspondence_S71 => state_S71, correspondence_C67 => state_C67, correspondence_S84 => state_S84, Sw03_state => state_Sw03, D04_state => state_D04, indication => signals_i(74), command => signals_o(74), correspondence_C125 => state_C125, clock => clock, reset => reset);
	railwaySignal_J38 : railwaySignal_75 port map(R23_command => cmd_R23_J38, R21_command => cmd_R21_J38, R87_command => cmd_R87_J38, track_ne996 => tracks_i(45), track_ne98 => tracks_i(20), correspondence_L30 => state_L30, correspondence_X50 => state_X50, indication => signals_i(75), command => signals_o(75), correspondence_J38 => state_J38, clock => clock, reset => reset);
	railwaySignal_S129 : railwaySignal_76 port map(R88_command => cmd_R88_S129, R89_command => cmd_R89_S129, R31_command => cmd_R31_S129, track_ne996 => tracks_i(45), track_ne292 => tracks_i(9), track_ne997 => tracks_i(46), track_ne297 => tracks_i(11), track_ne290 => tracks_i(8), track_ne384 => tracks_i(13), track_ne295 => tracks_i(10), correspondence_J37 => state_J37, correspondence_S71 => state_S71, correspondence_J35 => state_J35, correspondence_C67 => state_C67, correspondence_S84 => state_S84, Sw04_state => state_Sw04, D14_state => state_D14, Sw03_state => state_Sw03, D04_state => state_D04, indication => signals_i(76), command => signals_o(76), correspondence_S129 => state_S129, clock => clock, reset => reset);
	node_ne991 : node_0 port map(track_i => tracks_i(0), track_o => state_ne991, R1_command => cmd_R1_ne991, R20_command => cmd_R20_ne991, R39_command => cmd_R39_ne991, R40_command => cmd_R40_ne991, R41_command => cmd_R41_ne991, R60_command => cmd_R60_ne991, reset => reset);
	node_ne61 : node_1 port map(track_i => tracks_i(1), track_o => state_ne61, R35_command => cmd_R35_ne61, R51_command => cmd_R51_ne61, R53_command => cmd_R53_ne61, R54_command => cmd_R54_ne61, R64_command => cmd_R64_ne61, reset => reset);
	node_ne63 : node_2 port map(track_i => tracks_i(2), track_o => state_ne63, R4_command => cmd_R4_ne63, R34_command => cmd_R34_ne63, R36_command => cmd_R36_ne63, R65_command => cmd_R65_ne63, R66_command => cmd_R66_ne63, R67_command => cmd_R67_ne63, reset => reset);
	node_ne65 : node_3 port map(track_i => tracks_i(3), track_o => state_ne65, R65_command => cmd_R65_ne65, R66_command => cmd_R66_ne65, R79_command => cmd_R79_ne65, R80_command => cmd_R80_ne65, reset => reset);
	node_ne910 : node_4 port map(track_i => tracks_i(4), track_o => state_ne910, R38_command => cmd_R38_ne910, R55_command => cmd_R55_ne910, R57_command => cmd_R57_ne910, R58_command => cmd_R58_ne910, R77_command => cmd_R77_ne910, reset => reset);
	node_ne912 : node_5 port map(track_i => tracks_i(5), track_o => state_ne912, R8_command => cmd_R8_ne912, R26_command => cmd_R26_ne912, R28_command => cmd_R28_ne912, R37_command => cmd_R37_ne912, R75_command => cmd_R75_ne912, R76_command => cmd_R76_ne912, reset => reset);
	node_ne114 : node_6 port map(track_i => tracks_i(6), track_o => state_ne114, R10_command => cmd_R10_ne114, R17_command => cmd_R17_ne114, R27_command => cmd_R27_ne114, R29_command => cmd_R29_ne114, R68_command => cmd_R68_ne114, R69_command => cmd_R69_ne114, R70_command => cmd_R70_ne114, R71_command => cmd_R71_ne114, R73_command => cmd_R73_ne114, reset => reset);
	node_ne288 : node_7 port map(track_i => tracks_i(7), track_o => state_ne288, R39_command => cmd_R39_ne288, R41_command => cmd_R41_ne288, R43_command => cmd_R43_ne288, R44_command => cmd_R44_ne288, R60_command => cmd_R60_ne288, reset => reset);
	node_ne290 : node_8 port map(track_i => tracks_i(8), track_o => state_ne290, R2_command => cmd_R2_ne290, R20_command => cmd_R20_ne290, R22_command => cmd_R22_ne290, R40_command => cmd_R40_ne290, R61_command => cmd_R61_ne290, R62_command => cmd_R62_ne290, reset => reset);
	node_ne292 : node_9 port map(track_i => tracks_i(9), track_o => state_ne292, R21_command => cmd_R21_ne292, R22_command => cmd_R22_ne292, R61_command => cmd_R61_ne292, R88_command => cmd_R88_ne292, reset => reset);
	node_ne295 : node_10 port map(track_i => tracks_i(10), track_o => state_ne295, R41_command => cmd_R41_ne295, R43_command => cmd_R43_ne295, R45_command => cmd_R45_ne295, R46_command => cmd_R46_ne295, reset => reset);
	node_ne297 : node_11 port map(track_i => tracks_i(11), track_o => state_ne297, R11_command => cmd_R11_ne297, R42_command => cmd_R42_ne297, R45_command => cmd_R45_ne297, R46_command => cmd_R46_ne297, R47_command => cmd_R47_ne297, R85_command => cmd_R85_ne297, R86_command => cmd_R86_ne297, R87_command => cmd_R87_ne297, R89_command => cmd_R89_ne297, reset => reset);
	node_ne377 : node_12 port map(track_i => tracks_i(12), track_o => state_ne377, R2_command => cmd_R2_ne377, R3_command => cmd_R3_ne377, R12_command => cmd_R12_ne377, R62_command => cmd_R62_ne377, reset => reset);
	node_ne384 : node_13 port map(track_i => tracks_i(13), track_o => state_ne384, R11_command => cmd_R11_ne384, R42_command => cmd_R42_ne384, R47_command => cmd_R47_ne384, R59_command => cmd_R59_ne384, R60_command => cmd_R60_ne384, reset => reset);
	node_ne400 : node_14 port map(track_i => tracks_i(14), track_o => state_ne400, R13_command => cmd_R13_ne400, R48_command => cmd_R48_ne400, R49_command => cmd_R49_ne400, R50_command => cmd_R50_ne400, R52_command => cmd_R52_ne400, R81_command => cmd_R81_ne400, R82_command => cmd_R82_ne400, R83_command => cmd_R83_ne400, R84_command => cmd_R84_ne400, reset => reset);
	node_ne404 : node_15 port map(track_i => tracks_i(15), track_o => state_ne404, R48_command => cmd_R48_ne404, R49_command => cmd_R49_ne404, R51_command => cmd_R51_ne404, R53_command => cmd_R53_ne404, reset => reset);
	node_ne407 : node_16 port map(track_i => tracks_i(16), track_o => state_ne407, R13_command => cmd_R13_ne407, R50_command => cmd_R50_ne407, R52_command => cmd_R52_ne407, R63_command => cmd_R63_ne407, R64_command => cmd_R64_ne407, reset => reset);
	node_ne421 : node_17 port map(track_i => tracks_i(17), track_o => state_ne421, R4_command => cmd_R4_ne421, R5_command => cmd_R5_ne421, R14_command => cmd_R14_ne421, R67_command => cmd_R67_ne421, reset => reset);
	node_ne450 : node_18 port map(track_i => tracks_i(18), track_o => state_ne450, R6_command => cmd_R6_ne450, R7_command => cmd_R7_ne450, R72_command => cmd_R72_ne450, R74_command => cmd_R74_ne450, reset => reset);
	node_ne465 : node_19 port map(track_i => tracks_i(19), track_o => state_ne465, R8_command => cmd_R8_ne465, R9_command => cmd_R9_ne465, R15_command => cmd_R15_ne465, R75_command => cmd_R75_ne465, reset => reset);
	node_ne98 : node_20 port map(track_i => tracks_i(20), track_o => state_ne98, R18_command => cmd_R18_ne98, R23_command => cmd_R23_ne98, R30_command => cmd_R30_ne98, R31_command => cmd_R31_ne98, R34_command => cmd_R34_ne98, R51_command => cmd_R51_ne98, R64_command => cmd_R64_ne98, reset => reset);
	node_ne99 : node_21 port map(track_i => tracks_i(21), track_o => state_ne99, R30_command => cmd_R30_ne99, R34_command => cmd_R34_ne99, R35_command => cmd_R35_ne99, R36_command => cmd_R36_ne99, R51_command => cmd_R51_ne99, R64_command => cmd_R64_ne99, reset => reset);
	node_ne100 : node_22 port map(track_i => tracks_i(22), track_o => state_ne100, R19_command => cmd_R19_ne100, R24_command => cmd_R24_ne100, R25_command => cmd_R25_ne100, R32_command => cmd_R32_ne100, R33_command => cmd_R33_ne100, reset => reset);
	node_ne101 : node_23 port map(track_i => tracks_i(23), track_o => state_ne101, R25_command => cmd_R25_ne101, R26_command => cmd_R26_ne101, R32_command => cmd_R32_ne101, R37_command => cmd_R37_ne101, R38_command => cmd_R38_ne101, R55_command => cmd_R55_ne101, R77_command => cmd_R77_ne101, reset => reset);
	node_ne102 : node_24 port map(track_i => tracks_i(24), track_o => state_ne102, R10_command => cmd_R10_ne102, R29_command => cmd_R29_ne102, reset => reset);
	node_ne104 : node_25 port map(track_i => tracks_i(25), track_o => state_ne104, R11_command => cmd_R11_ne104, R59_command => cmd_R59_ne104, reset => reset);
	node_ne110 : node_26 port map(track_i => tracks_i(26), track_o => state_ne110, R42_command => cmd_R42_ne110, R44_command => cmd_R44_ne110, R60_command => cmd_R60_ne110, reset => reset);
	node_ne111 : node_27 port map(track_i => tracks_i(27), track_o => state_ne111, R2_command => cmd_R2_ne111, R62_command => cmd_R62_ne111, reset => reset);
	node_ne113 : node_28 port map(track_i => tracks_i(28), track_o => state_ne113, R3_command => cmd_R3_ne113, R12_command => cmd_R12_ne113, reset => reset);
	node_ne122 : node_29 port map(track_i => tracks_i(29), track_o => state_ne122, R13_command => cmd_R13_ne122, R63_command => cmd_R63_ne122, reset => reset);
	node_ne123 : node_30 port map(track_i => tracks_i(30), track_o => state_ne123, R52_command => cmd_R52_ne123, R54_command => cmd_R54_ne123, R64_command => cmd_R64_ne123, reset => reset);
	node_ne124 : node_31 port map(track_i => tracks_i(31), track_o => state_ne124, R4_command => cmd_R4_ne124, R67_command => cmd_R67_ne124, reset => reset);
	node_ne126 : node_32 port map(track_i => tracks_i(32), track_o => state_ne126, R5_command => cmd_R5_ne126, R14_command => cmd_R14_ne126, reset => reset);
	node_ne127 : node_33 port map(track_i => tracks_i(33), track_o => state_ne127, R6_command => cmd_R6_ne127, R16_command => cmd_R16_ne127, R56_command => cmd_R56_ne127, R69_command => cmd_R69_ne127, R71_command => cmd_R71_ne127, R72_command => cmd_R72_ne127, R77_command => cmd_R77_ne127, R78_command => cmd_R78_ne127, reset => reset);
	node_ne129 : node_34 port map(track_i => tracks_i(34), track_o => state_ne129, R69_command => cmd_R69_ne129, R70_command => cmd_R70_ne129, R71_command => cmd_R71_ne129, R73_command => cmd_R73_ne129, reset => reset);
	node_ne130 : node_35 port map(track_i => tracks_i(35), track_o => state_ne130, R7_command => cmd_R7_ne130, R55_command => cmd_R55_ne130, R57_command => cmd_R57_ne130, R70_command => cmd_R70_ne130, R73_command => cmd_R73_ne130, R74_command => cmd_R74_ne130, reset => reset);
	node_ne131 : node_36 port map(track_i => tracks_i(36), track_o => state_ne131, R8_command => cmd_R8_ne131, R75_command => cmd_R75_ne131, reset => reset);
	node_ne132 : node_37 port map(track_i => tracks_i(37), track_o => state_ne132, R27_command => cmd_R27_ne132, R28_command => cmd_R28_ne132, R68_command => cmd_R68_ne132, R76_command => cmd_R76_ne132, reset => reset);
	node_ne133 : node_38 port map(track_i => tracks_i(38), track_o => state_ne133, R9_command => cmd_R9_ne133, R15_command => cmd_R15_ne133, reset => reset);
	node_ne134 : node_39 port map(track_i => tracks_i(39), track_o => state_ne134, R16_command => cmd_R16_ne134, R78_command => cmd_R78_ne134, reset => reset);
	node_ne135 : node_40 port map(track_i => tracks_i(40), track_o => state_ne135, R56_command => cmd_R56_ne135, R58_command => cmd_R58_ne135, R77_command => cmd_R77_ne135, reset => reset);
	node_ne992 : node_41 port map(track_i => tracks_i(41), track_o => state_ne992, R24_command => cmd_R24_ne992, R33_command => cmd_R33_ne992, R79_command => cmd_R79_ne992, R80_command => cmd_R80_ne992, R81_command => cmd_R81_ne992, R84_command => cmd_R84_ne992, reset => reset);
	node_ne993 : node_42 port map(track_i => tracks_i(42), track_o => state_ne993, R82_command => cmd_R82_ne993, R83_command => cmd_R83_ne993, reset => reset);
	node_ne994 : node_43 port map(track_i => tracks_i(43), track_o => state_ne994, R81_command => cmd_R81_ne994, R84_command => cmd_R84_ne994, reset => reset);
	node_ne995 : node_44 port map(track_i => tracks_i(44), track_o => state_ne995, R85_command => cmd_R85_ne995, R86_command => cmd_R86_ne995, reset => reset);
	node_ne996 : node_45 port map(track_i => tracks_i(45), track_o => state_ne996, R21_command => cmd_R21_ne996, R23_command => cmd_R23_ne996, R31_command => cmd_R31_ne996, R87_command => cmd_R87_ne996, R88_command => cmd_R88_ne996, R89_command => cmd_R89_ne996, reset => reset);
	node_ne997 : node_46 port map(track_i => tracks_i(46), track_o => state_ne997, R87_command => cmd_R87_ne997, R89_command => cmd_R89_ne997, reset => reset);
	route_R1 : route_0 port map(routeRequest => routes_i(0), ne991_command => cmd_R1_ne991, track_ne991 => state_ne991, D01_command => cmd_R1_D01, D01_state => state_D01, T02_state => state_T02, T02_command => cmd_R1_T02, S64_state => state_S64, S64_command =>cmd_R1_S64, routeExecute => routes_o(0), clock => clock, reset => reset);
	route_R2 : route_1 port map(routeRequest => routes_i(1), ne290_command => cmd_R2_ne290, track_ne290 => state_ne290, ne377_command => cmd_R2_ne377, track_ne377 => state_ne377, ne111_command => cmd_R2_ne111, track_ne111 => state_ne111, D01_command => cmd_R2_D01, D01_state => state_D01, D14_command => cmd_R2_D14, D14_state => state_D14, D15_command => cmd_R2_D15, D15_state => state_D15, T04_state => state_T04, T04_command => cmd_R2_T04, J35_state => state_J35, J35_command =>cmd_R2_J35, routeExecute => routes_o(1), clock => clock, reset => reset);
	route_R3 : route_2 port map(routeRequest => routes_i(2), ne377_command => cmd_R3_ne377, track_ne377 => state_ne377, ne113_command => cmd_R3_ne113, track_ne113 => state_ne113, D15_command => cmd_R3_D15, D15_state => state_D15, T04_state => state_T04, T04_command => cmd_R3_T04, T15_state => state_T15, T15_command =>cmd_R3_T15, routeExecute => routes_o(2), clock => clock, reset => reset);
	route_R4 : route_3 port map(routeRequest => routes_i(3), ne63_command => cmd_R4_ne63, track_ne63 => state_ne63, ne421_command => cmd_R4_ne421, track_ne421 => state_ne421, ne124_command => cmd_R4_ne124, track_ne124 => state_ne124, D05_command => cmd_R4_D05, D05_state => state_D05, D18_command => cmd_R4_D18, D18_state => state_D18, D19_command => cmd_R4_D19, D19_state => state_D19, T06_state => state_T06, T06_command => cmd_R4_T06, C54_state => state_C54, C54_command =>cmd_R4_C54, routeExecute => routes_o(3), clock => clock, reset => reset);
	route_R5 : route_4 port map(routeRequest => routes_i(4), ne421_command => cmd_R5_ne421, track_ne421 => state_ne421, ne126_command => cmd_R5_ne126, track_ne126 => state_ne126, D19_command => cmd_R5_D19, D19_state => state_D19, T06_state => state_T06, T06_command => cmd_R5_T06, T19_state => state_T19, T19_command =>cmd_R5_T19, routeExecute => routes_o(4), clock => clock, reset => reset);
	route_R6 : route_5 port map(routeRequest => routes_i(5), ne450_command => cmd_R6_ne450, track_ne450 => state_ne450, ne127_command => cmd_R6_ne127, track_ne127 => state_ne127, D10_command => cmd_R6_D10, D10_state => state_D10, D09_command => cmd_R6_D09, D09_state => state_D09, D24_command => cmd_R6_D24, D24_state => state_D24, D12_command => cmd_R6_D12, D12_state => state_D12, T08_state => state_T08, T08_command => cmd_R6_T08, S117_state => state_S117, S117_command =>cmd_R6_S117, routeExecute => routes_o(5), clock => clock, reset => reset);
	route_R7 : route_6 port map(routeRequest => routes_i(6), ne450_command => cmd_R7_ne450, track_ne450 => state_ne450, ne130_command => cmd_R7_ne130, track_ne130 => state_ne130, D10_command => cmd_R7_D10, D10_state => state_D10, D09_command => cmd_R7_D09, D09_state => state_D09, D12_command => cmd_R7_D12, D12_state => state_D12, T08_state => state_T08, T08_command => cmd_R7_T08, C79_state => state_C79, C79_command =>cmd_R7_C79, routeExecute => routes_o(6), clock => clock, reset => reset);
	route_R8 : route_7 port map(routeRequest => routes_i(7), ne912_command => cmd_R8_ne912, track_ne912 => state_ne912, ne465_command => cmd_R8_ne465, track_ne465 => state_ne465, ne131_command => cmd_R8_ne131, track_ne131 => state_ne131, D09_command => cmd_R8_D09, D09_state => state_D09, D20_command => cmd_R8_D20, D20_state => state_D20, D21_command => cmd_R8_D21, D21_state => state_D21, T10_state => state_T10, T10_command => cmd_R8_T10, J45_state => state_J45, J45_command =>cmd_R8_J45, routeExecute => routes_o(7), clock => clock, reset => reset);
	route_R9 : route_8 port map(routeRequest => routes_i(8), ne465_command => cmd_R9_ne465, track_ne465 => state_ne465, ne133_command => cmd_R9_ne133, track_ne133 => state_ne133, D21_command => cmd_R9_D21, D21_state => state_D21, T10_state => state_T10, T10_command => cmd_R9_T10, T21_state => state_T21, T21_command =>cmd_R9_T21, routeExecute => routes_o(8), clock => clock, reset => reset);
	route_R10 : route_9 port map(routeRequest => routes_i(9), ne114_command => cmd_R10_ne114, track_ne114 => state_ne114, ne102_command => cmd_R10_ne102, track_ne102 => state_ne102, D23_command => cmd_R10_D23, D23_state => state_D23, T12_state => state_T12, T12_command => cmd_R10_T12, S101_state => state_S101, S101_command =>cmd_R10_S101, routeExecute => routes_o(9), clock => clock, reset => reset);
	route_R11 : route_10 port map(routeRequest => routes_i(10), ne297_command => cmd_R11_ne297, track_ne297 => state_ne297, ne384_command => cmd_R11_ne384, track_ne384 => state_ne384, ne104_command => cmd_R11_ne104, track_ne104 => state_ne104, D04_command => cmd_R11_D04, D04_state => state_D04, Sw03_command => cmd_R11_Sw03, Sw03_state => state_Sw03, Sw02_command => cmd_R11_Sw02, Sw02_state => state_Sw02, T14_state => state_T14, T14_command => cmd_R11_T14, S126_state => state_S126, S126_command =>cmd_R11_S126, routeExecute => routes_o(10), clock => clock, reset => reset);
	route_R12 : route_11 port map(routeRequest => routes_i(11), ne377_command => cmd_R12_ne377, track_ne377 => state_ne377, ne113_command => cmd_R12_ne113, track_ne113 => state_ne113, D15_command => cmd_R12_D15, D15_state => state_D15, T16_state => state_T16, T16_command => cmd_R12_T16, T03_state => state_T03, T03_command =>cmd_R12_T03, routeExecute => routes_o(11), clock => clock, reset => reset);
	route_R13 : route_12 port map(routeRequest => routes_i(12), ne400_command => cmd_R13_ne400, track_ne400 => state_ne400, ne407_command => cmd_R13_ne407, track_ne407 => state_ne407, ne122_command => cmd_R13_ne122, track_ne122 => state_ne122, D07_command => cmd_R13_D07, D07_state => state_D07, Sw05_command => cmd_R13_Sw05, Sw05_state => state_Sw05, D16_command => cmd_R13_D16, D16_state => state_D16, T18_state => state_T18, T18_command => cmd_R13_T18, S123_state => state_S123, S123_command =>cmd_R13_S123, routeExecute => routes_o(12), clock => clock, reset => reset);
	route_R14 : route_13 port map(routeRequest => routes_i(13), ne421_command => cmd_R14_ne421, track_ne421 => state_ne421, ne126_command => cmd_R14_ne126, track_ne126 => state_ne126, D19_command => cmd_R14_D19, D19_state => state_D19, T20_state => state_T20, T20_command => cmd_R14_T20, T05_state => state_T05, T05_command =>cmd_R14_T05, routeExecute => routes_o(13), clock => clock, reset => reset);
	route_R15 : route_14 port map(routeRequest => routes_i(14), ne465_command => cmd_R15_ne465, track_ne465 => state_ne465, ne133_command => cmd_R15_ne133, track_ne133 => state_ne133, D21_command => cmd_R15_D21, D21_state => state_D21, T22_state => state_T22, T22_command => cmd_R15_T22, T09_state => state_T09, T09_command =>cmd_R15_T09, routeExecute => routes_o(14), clock => clock, reset => reset);
	route_R16 : route_15 port map(routeRequest => routes_i(15), ne127_command => cmd_R16_ne127, track_ne127 => state_ne127, ne134_command => cmd_R16_ne134, track_ne134 => state_ne134, D23_command => cmd_R16_D23, D23_state => state_D23, D24_command => cmd_R16_D24, D24_state => state_D24, T24_state => state_T24, T24_command => cmd_R16_T24, S104_state => state_S104, S104_command =>cmd_R16_S104, routeExecute => routes_o(15), clock => clock, reset => reset);
	route_R17 : route_16 port map(routeRequest => routes_i(16), ne114_command => cmd_R17_ne114, track_ne114 => state_ne114, L29_state => state_L29, L29_command => cmd_R17_L29, J48_state => state_J48, J48_command =>cmd_R17_J48, routeExecute => routes_o(16), clock => clock, reset => reset);
	route_R18 : route_17 port map(routeRequest => routes_i(17), ne98_command => cmd_R18_ne98, track_ne98 => state_ne98, L30_state => state_L30, L30_command => cmd_R18_L30, X50_state => state_X50, X50_command =>cmd_R18_X50, routeExecute => routes_o(17), clock => clock, reset => reset);
	route_R19 : route_18 port map(routeRequest => routes_i(18), ne100_command => cmd_R19_ne100, track_ne100 => state_ne100, L31_state => state_L31, L31_command => cmd_R19_L31, X52_state => state_X52, X52_command =>cmd_R19_X52, routeExecute => routes_o(18), clock => clock, reset => reset);
	route_R20 : route_19 port map(routeRequest => routes_i(19), ne991_command => cmd_R20_ne991, track_ne991 => state_ne991, ne290_command => cmd_R20_ne290, track_ne290 => state_ne290, D01_command => cmd_R20_D01, D01_state => state_D01, J35_state => state_J35, J35_command => cmd_R20_J35, T01_state => state_T01, T01_command =>cmd_R20_T01, routeExecute => routes_o(19), clock => clock, reset => reset);
	route_R21 : route_20 port map(routeRequest => routes_i(20), ne292_command => cmd_R21_ne292, track_ne292 => state_ne292, ne996_command => cmd_R21_ne996, track_ne996 => state_ne996, Sw04_command => cmd_R21_Sw04, Sw04_state => state_Sw04, J36_state => state_J36, J36_command => cmd_R21_J36, J38_state => state_J38, J38_command =>cmd_R21_J38, routeExecute => routes_o(20), clock => clock, reset => reset);
	route_R22 : route_21 port map(routeRequest => routes_i(21), ne290_command => cmd_R22_ne290, track_ne290 => state_ne290, ne292_command => cmd_R22_ne292, track_ne292 => state_ne292, D01_command => cmd_R22_D01, D01_state => state_D01, D14_command => cmd_R22_D14, D14_state => state_D14, J37_state => state_J37, J37_command => cmd_R22_J37, J35_state => state_J35, J35_command =>cmd_R22_J35, routeExecute => routes_o(21), clock => clock, reset => reset);
	route_R23 : route_22 port map(routeRequest => routes_i(22), ne98_command => cmd_R23_ne98, track_ne98 => state_ne98, ne996_command => cmd_R23_ne996, track_ne996 => state_ne996, J38_state => state_J38, J38_command => cmd_R23_J38, L30_state => state_L30, L30_command =>cmd_R23_L30, routeExecute => routes_o(22), clock => clock, reset => reset);
	route_R24 : route_23 port map(routeRequest => routes_i(23), ne100_command => cmd_R24_ne100, track_ne100 => state_ne100, ne992_command => cmd_R24_ne992, track_ne992 => state_ne992, J40_state => state_J40, J40_command => cmd_R24_J40, L31_state => state_L31, L31_command =>cmd_R24_L31, routeExecute => routes_o(23), clock => clock, reset => reset);
	route_R25 : route_24 port map(routeRequest => routes_i(24), ne100_command => cmd_R25_ne100, track_ne100 => state_ne100, ne101_command => cmd_R25_ne101, track_ne101 => state_ne101, J43_state => state_J43, J43_command => cmd_R25_J43, X53_state => state_X53, X53_command =>cmd_R25_X53, routeExecute => routes_o(24), clock => clock, reset => reset);
	route_R26 : route_25 port map(routeRequest => routes_i(25), ne912_command => cmd_R26_ne912, track_ne912 => state_ne912, ne101_command => cmd_R26_ne101, track_ne101 => state_ne101, D09_command => cmd_R26_D09, D09_state => state_D09, J45_state => state_J45, J45_command => cmd_R26_J45, J43_state => state_J43, J43_command =>cmd_R26_J43, routeExecute => routes_o(25), clock => clock, reset => reset);
	route_R27 : route_26 port map(routeRequest => routes_i(26), ne114_command => cmd_R27_ne114, track_ne114 => state_ne114, ne132_command => cmd_R27_ne132, track_ne132 => state_ne132, D23_command => cmd_R27_D23, D23_state => state_D23, J46_state => state_J46, J46_command => cmd_R27_J46, L29_state => state_L29, L29_command =>cmd_R27_L29, routeExecute => routes_o(26), clock => clock, reset => reset);
	route_R28 : route_27 port map(routeRequest => routes_i(27), ne912_command => cmd_R28_ne912, track_ne912 => state_ne912, ne132_command => cmd_R28_ne132, track_ne132 => state_ne132, D09_command => cmd_R28_D09, D09_state => state_D09, D20_command => cmd_R28_D20, D20_state => state_D20, J47_state => state_J47, J47_command => cmd_R28_J47, J45_state => state_J45, J45_command =>cmd_R28_J45, routeExecute => routes_o(27), clock => clock, reset => reset);
	route_R29 : route_28 port map(routeRequest => routes_i(28), ne114_command => cmd_R29_ne114, track_ne114 => state_ne114, ne102_command => cmd_R29_ne102, track_ne102 => state_ne102, J48_state => state_J48, J48_command => cmd_R29_J48, T11_state => state_T11, T11_command =>cmd_R29_T11, routeExecute => routes_o(28), clock => clock, reset => reset);
	route_R30 : route_29 port map(routeRequest => routes_i(29), ne98_command => cmd_R30_ne98, track_ne98 => state_ne98, ne99_command => cmd_R30_ne99, track_ne99 => state_ne99, Lc01_command => cmd_R30_Lc01, Lc01_state => state_Lc01, D05_command => cmd_R30_D05, D05_state => state_D05, X50_state => state_X50, X50_command => cmd_R30_X50, S55_state => state_S55, S55_command =>cmd_R30_S55, routeExecute => routes_o(29), clock => clock, reset => reset);
	route_R31 : route_30 port map(routeRequest => routes_i(30), ne98_command => cmd_R31_ne98, track_ne98 => state_ne98, ne996_command => cmd_R31_ne996, track_ne996 => state_ne996, Lc01_command => cmd_R31_Lc01, Lc01_state => state_Lc01, Sw04_command => cmd_R31_Sw04, Sw04_state => state_Sw04, Sw03_command => cmd_R31_Sw03, Sw03_state => state_Sw03, X51_state => state_X51, X51_command => cmd_R31_X51, S129_state => state_S129, S129_command =>cmd_R31_S129, routeExecute => routes_o(30), clock => clock, reset => reset);
	route_R32 : route_31 port map(routeRequest => routes_i(31), ne100_command => cmd_R32_ne100, track_ne100 => state_ne100, ne101_command => cmd_R32_ne101, track_ne101 => state_ne101, Lc04_command => cmd_R32_Lc04, Lc04_state => state_Lc04, D09_command => cmd_R32_D09, D09_state => state_D09, X52_state => state_X52, X52_command => cmd_R32_X52, S59_state => state_S59, S59_command =>cmd_R32_S59, routeExecute => routes_o(31), clock => clock, reset => reset);
	route_R33 : route_32 port map(routeRequest => routes_i(32), ne100_command => cmd_R33_ne100, track_ne100 => state_ne100, ne992_command => cmd_R33_ne992, track_ne992 => state_ne992, Lc04_command => cmd_R33_Lc04, Lc04_state => state_Lc04, Sw01_command => cmd_R33_Sw01, Sw01_state => state_Sw01, Sw05_command => cmd_R33_Sw05, Sw05_state => state_Sw05, X53_state => state_X53, X53_command => cmd_R33_X53, S120_state => state_S120, S120_command =>cmd_R33_S120, routeExecute => routes_o(32), clock => clock, reset => reset);
	route_R34 : route_33 port map(routeRequest => routes_i(33), ne63_command => cmd_R34_ne63, track_ne63 => state_ne63, ne98_command => cmd_R34_ne98, track_ne98 => state_ne98, ne99_command => cmd_R34_ne99, track_ne99 => state_ne99, Lc01_command => cmd_R34_Lc01, Lc01_state => state_Lc01, D05_command => cmd_R34_D05, D05_state => state_D05, C54_state => state_C54, C54_command => cmd_R34_C54, X51_state => state_X51, X51_command =>cmd_R34_X51, routeExecute => routes_o(33), clock => clock, reset => reset);
	route_R35 : route_34 port map(routeRequest => routes_i(34), ne61_command => cmd_R35_ne61, track_ne61 => state_ne61, ne99_command => cmd_R35_ne99, track_ne99 => state_ne99, D08_command => cmd_R35_D08, D08_state => state_D08, D05_command => cmd_R35_D05, D05_state => state_D05, S55_state => state_S55, S55_command => cmd_R35_S55, S78_state => state_S78, S78_command =>cmd_R35_S78, routeExecute => routes_o(34), clock => clock, reset => reset);
	route_R36 : route_35 port map(routeRequest => routes_i(35), ne63_command => cmd_R36_ne63, track_ne63 => state_ne63, ne99_command => cmd_R36_ne99, track_ne99 => state_ne99, D05_command => cmd_R36_D05, D05_state => state_D05, D18_command => cmd_R36_D18, D18_state => state_D18, S55_state => state_S55, S55_command => cmd_R36_S55, S95_state => state_S95, S95_command =>cmd_R36_S95, routeExecute => routes_o(35), clock => clock, reset => reset);
	route_R37 : route_36 port map(routeRequest => routes_i(36), ne912_command => cmd_R37_ne912, track_ne912 => state_ne912, ne101_command => cmd_R37_ne101, track_ne101 => state_ne101, D09_command => cmd_R37_D09, D09_state => state_D09, D20_command => cmd_R37_D20, D20_state => state_D20, D21_command => cmd_R37_D21, D21_state => state_D21, S59_state => state_S59, S59_command => cmd_R37_S59, S110_state => state_S110, S110_command =>cmd_R37_S110, routeExecute => routes_o(36), clock => clock, reset => reset);
	route_R38 : route_37 port map(routeRequest => routes_i(37), ne910_command => cmd_R38_ne910, track_ne910 => state_ne910, ne101_command => cmd_R38_ne101, track_ne101 => state_ne101, D10_command => cmd_R38_D10, D10_state => state_D10, D09_command => cmd_R38_D09, D09_state => state_D09, S59_state => state_S59, S59_command => cmd_R38_S59, S81_state => state_S81, S81_command =>cmd_R38_S81, routeExecute => routes_o(37), clock => clock, reset => reset);
	route_R39 : route_38 port map(routeRequest => routes_i(38), ne991_command => cmd_R39_ne991, track_ne991 => state_ne991, ne288_command => cmd_R39_ne288, track_ne288 => state_ne288, D01_command => cmd_R39_D01, D01_state => state_D01, D03_command => cmd_R39_D03, D03_state => state_D03, S64_state => state_S64, S64_command => cmd_R39_S64, S69_state => state_S69, S69_command =>cmd_R39_S69, routeExecute => routes_o(38), clock => clock, reset => reset);
	route_R40 : route_39 port map(routeRequest => routes_i(39), ne991_command => cmd_R40_ne991, track_ne991 => state_ne991, ne290_command => cmd_R40_ne290, track_ne290 => state_ne290, D01_command => cmd_R40_D01, D01_state => state_D01, D14_command => cmd_R40_D14, D14_state => state_D14, S64_state => state_S64, S64_command => cmd_R40_S64, S86_state => state_S86, S86_command =>cmd_R40_S86, routeExecute => routes_o(39), clock => clock, reset => reset);
	route_R41 : route_40 port map(routeRequest => routes_i(40), ne991_command => cmd_R41_ne991, track_ne991 => state_ne991, ne288_command => cmd_R41_ne288, track_ne288 => state_ne288, ne295_command => cmd_R41_ne295, track_ne295 => state_ne295, D01_command => cmd_R41_D01, D01_state => state_D01, D03_command => cmd_R41_D03, D03_state => state_D03, C67_state => state_C67, C67_command => cmd_R41_C67, T01_state => state_T01, T01_command =>cmd_R41_T01, routeExecute => routes_o(40), clock => clock, reset => reset);
	route_R42 : route_41 port map(routeRequest => routes_i(41), ne297_command => cmd_R42_ne297, track_ne297 => state_ne297, ne384_command => cmd_R42_ne384, track_ne384 => state_ne384, ne110_command => cmd_R42_ne110, track_ne110 => state_ne110, D04_command => cmd_R42_D04, D04_state => state_D04, Sw03_command => cmd_R42_Sw03, Sw03_state => state_Sw03, Sw02_command => cmd_R42_Sw02, Sw02_state => state_Sw02, B68_state => state_B68, B68_command => cmd_R42_B68, S126_state => state_S126, S126_command =>cmd_R42_S126, routeExecute => routes_o(41), clock => clock, reset => reset);
	route_R43 : route_42 port map(routeRequest => routes_i(42), ne288_command => cmd_R43_ne288, track_ne288 => state_ne288, ne295_command => cmd_R43_ne295, track_ne295 => state_ne295, D03_command => cmd_R43_D03, D03_state => state_D03, D04_command => cmd_R43_D04, D04_state => state_D04, S69_state => state_S69, S69_command => cmd_R43_S69, C70_state => state_C70, C70_command =>cmd_R43_C70, routeExecute => routes_o(42), clock => clock, reset => reset);
	route_R44 : route_43 port map(routeRequest => routes_i(43), ne288_command => cmd_R44_ne288, track_ne288 => state_ne288, ne110_command => cmd_R44_ne110, track_ne110 => state_ne110, D03_command => cmd_R44_D03, D03_state => state_D03, D04_command => cmd_R44_D04, D04_state => state_D04, Sw02_command => cmd_R44_Sw02, Sw02_state => state_Sw02, S69_state => state_S69, S69_command => cmd_R44_S69, B68_state => state_B68, B68_command =>cmd_R44_B68, routeExecute => routes_o(43), clock => clock, reset => reset);
	route_R45 : route_44 port map(routeRequest => routes_i(44), ne295_command => cmd_R45_ne295, track_ne295 => state_ne295, ne297_command => cmd_R45_ne297, track_ne297 => state_ne297, D04_command => cmd_R45_D04, D04_state => state_D04, Sw03_command => cmd_R45_Sw03, Sw03_state => state_Sw03, C70_state => state_C70, C70_command => cmd_R45_C70, S126_state => state_S126, S126_command =>cmd_R45_S126, routeExecute => routes_o(44), clock => clock, reset => reset);
	route_R46 : route_45 port map(routeRequest => routes_i(45), ne295_command => cmd_R46_ne295, track_ne295 => state_ne295, ne297_command => cmd_R46_ne297, track_ne297 => state_ne297, D01_command => cmd_R46_D01, D01_state => state_D01, D03_command => cmd_R46_D03, D03_state => state_D03, D04_command => cmd_R46_D04, D04_state => state_D04, S71_state => state_S71, S71_command => cmd_R46_S71, C67_state => state_C67, C67_command =>cmd_R46_C67, routeExecute => routes_o(45), clock => clock, reset => reset);
	route_R47 : route_46 port map(routeRequest => routes_i(46), ne297_command => cmd_R47_ne297, track_ne297 => state_ne297, ne384_command => cmd_R47_ne384, track_ne384 => state_ne384, D04_command => cmd_R47_D04, D04_state => state_D04, Sw02_command => cmd_R47_Sw02, Sw02_state => state_Sw02, S71_state => state_S71, S71_command => cmd_R47_S71, S84_state => state_S84, S84_command =>cmd_R47_S84, routeExecute => routes_o(46), clock => clock, reset => reset);
	route_R48 : route_47 port map(routeRequest => routes_i(47), ne400_command => cmd_R48_ne400, track_ne400 => state_ne400, ne404_command => cmd_R48_ne404, track_ne404 => state_ne404, D07_command => cmd_R48_D07, D07_state => state_D07, Sw05_command => cmd_R48_Sw05, Sw05_state => state_Sw05, C73_state => state_C73, C73_command => cmd_R48_C73, S123_state => state_S123, S123_command =>cmd_R48_S123, routeExecute => routes_o(47), clock => clock, reset => reset);
	route_R49 : route_48 port map(routeRequest => routes_i(48), ne400_command => cmd_R49_ne400, track_ne400 => state_ne400, ne404_command => cmd_R49_ne404, track_ne404 => state_ne404, D08_command => cmd_R49_D08, D08_state => state_D08, D05_command => cmd_R49_D05, D05_state => state_D05, D07_command => cmd_R49_D07, D07_state => state_D07, S74_state => state_S74, S74_command => cmd_R49_S74, C76_state => state_C76, C76_command =>cmd_R49_C76, routeExecute => routes_o(48), clock => clock, reset => reset);
	route_R50 : route_49 port map(routeRequest => routes_i(49), ne400_command => cmd_R50_ne400, track_ne400 => state_ne400, ne407_command => cmd_R50_ne407, track_ne407 => state_ne407, D07_command => cmd_R50_D07, D07_state => state_D07, D16_command => cmd_R50_D16, D16_state => state_D16, S74_state => state_S74, S74_command => cmd_R50_S74, S93_state => state_S93, S93_command =>cmd_R50_S93, routeExecute => routes_o(49), clock => clock, reset => reset);
	route_R51 : route_50 port map(routeRequest => routes_i(50), ne61_command => cmd_R51_ne61, track_ne61 => state_ne61, ne404_command => cmd_R51_ne404, track_ne404 => state_ne404, ne98_command => cmd_R51_ne98, track_ne98 => state_ne98, ne99_command => cmd_R51_ne99, track_ne99 => state_ne99, Lc01_command => cmd_R51_Lc01, Lc01_state => state_Lc01, D08_command => cmd_R51_D08, D08_state => state_D08, D05_command => cmd_R51_D05, D05_state => state_D05, C76_state => state_C76, C76_command => cmd_R51_C76, X51_state => state_X51, X51_command =>cmd_R51_X51, routeExecute => routes_o(50), clock => clock, reset => reset);
	route_R52 : route_51 port map(routeRequest => routes_i(51), ne400_command => cmd_R52_ne400, track_ne400 => state_ne400, ne407_command => cmd_R52_ne407, track_ne407 => state_ne407, ne123_command => cmd_R52_ne123, track_ne123 => state_ne123, D07_command => cmd_R52_D07, D07_state => state_D07, Sw05_command => cmd_R52_Sw05, Sw05_state => state_Sw05, D16_command => cmd_R52_D16, D16_state => state_D16, B77_state => state_B77, B77_command => cmd_R52_B77, S123_state => state_S123, S123_command =>cmd_R52_S123, routeExecute => routes_o(51), clock => clock, reset => reset);
	route_R53 : route_52 port map(routeRequest => routes_i(52), ne61_command => cmd_R53_ne61, track_ne61 => state_ne61, ne404_command => cmd_R53_ne404, track_ne404 => state_ne404, D08_command => cmd_R53_D08, D08_state => state_D08, D07_command => cmd_R53_D07, D07_state => state_D07, S78_state => state_S78, S78_command => cmd_R53_S78, C73_state => state_C73, C73_command =>cmd_R53_C73, routeExecute => routes_o(52), clock => clock, reset => reset);
	route_R54 : route_53 port map(routeRequest => routes_i(53), ne61_command => cmd_R54_ne61, track_ne61 => state_ne61, ne123_command => cmd_R54_ne123, track_ne123 => state_ne123, D08_command => cmd_R54_D08, D08_state => state_D08, D07_command => cmd_R54_D07, D07_state => state_D07, D16_command => cmd_R54_D16, D16_state => state_D16, S78_state => state_S78, S78_command => cmd_R54_S78, B77_state => state_B77, B77_command =>cmd_R54_B77, routeExecute => routes_o(53), clock => clock, reset => reset);
	route_R55 : route_54 port map(routeRequest => routes_i(54), ne910_command => cmd_R55_ne910, track_ne910 => state_ne910, ne101_command => cmd_R55_ne101, track_ne101 => state_ne101, ne130_command => cmd_R55_ne130, track_ne130 => state_ne130, D10_command => cmd_R55_D10, D10_state => state_D10, D09_command => cmd_R55_D09, D09_state => state_D09, C79_state => state_C79, C79_command => cmd_R55_C79, J43_state => state_J43, J43_command =>cmd_R55_J43, routeExecute => routes_o(54), clock => clock, reset => reset);
	route_R56 : route_55 port map(routeRequest => routes_i(55), ne127_command => cmd_R56_ne127, track_ne127 => state_ne127, ne135_command => cmd_R56_ne135, track_ne135 => state_ne135, D23_command => cmd_R56_D23, D23_state => state_D23, D24_command => cmd_R56_D24, D24_state => state_D24, B80_state => state_B80, B80_command => cmd_R56_B80, S104_state => state_S104, S104_command =>cmd_R56_S104, routeExecute => routes_o(55), clock => clock, reset => reset);
	route_R57 : route_56 port map(routeRequest => routes_i(56), ne910_command => cmd_R57_ne910, track_ne910 => state_ne910, ne130_command => cmd_R57_ne130, track_ne130 => state_ne130, D10_command => cmd_R57_D10, D10_state => state_D10, D23_command => cmd_R57_D23, D23_state => state_D23, S81_state => state_S81, S81_command => cmd_R57_S81, S107_state => state_S107, S107_command =>cmd_R57_S107, routeExecute => routes_o(56), clock => clock, reset => reset);
	route_R58 : route_57 port map(routeRequest => routes_i(57), ne910_command => cmd_R58_ne910, track_ne910 => state_ne910, ne135_command => cmd_R58_ne135, track_ne135 => state_ne135, D10_command => cmd_R58_D10, D10_state => state_D10, D24_command => cmd_R58_D24, D24_state => state_D24, S81_state => state_S81, S81_command => cmd_R58_S81, B80_state => state_B80, B80_command =>cmd_R58_B80, routeExecute => routes_o(57), clock => clock, reset => reset);
	route_R59 : route_58 port map(routeRequest => routes_i(58), ne384_command => cmd_R59_ne384, track_ne384 => state_ne384, ne104_command => cmd_R59_ne104, track_ne104 => state_ne104, Sw02_command => cmd_R59_Sw02, Sw02_state => state_Sw02, S84_state => state_S84, S84_command => cmd_R59_S84, T13_state => state_T13, T13_command =>cmd_R59_T13, routeExecute => routes_o(58), clock => clock, reset => reset);
	route_R60 : route_59 port map(routeRequest => routes_i(59), ne991_command => cmd_R60_ne991, track_ne991 => state_ne991, ne288_command => cmd_R60_ne288, track_ne288 => state_ne288, ne384_command => cmd_R60_ne384, track_ne384 => state_ne384, ne110_command => cmd_R60_ne110, track_ne110 => state_ne110, D01_command => cmd_R60_D01, D01_state => state_D01, D03_command => cmd_R60_D03, D03_state => state_D03, Sw02_command => cmd_R60_Sw02, Sw02_state => state_Sw02, S84_state => state_S84, S84_command => cmd_R60_S84, T01_state => state_T01, T01_command =>cmd_R60_T01, routeExecute => routes_o(59), clock => clock, reset => reset);
	route_R61 : route_60 port map(routeRequest => routes_i(60), ne290_command => cmd_R61_ne290, track_ne290 => state_ne290, ne292_command => cmd_R61_ne292, track_ne292 => state_ne292, D14_command => cmd_R61_D14, D14_state => state_D14, Sw04_command => cmd_R61_Sw04, Sw04_state => state_Sw04, S86_state => state_S86, S86_command => cmd_R61_S86, J36_state => state_J36, J36_command =>cmd_R61_J36, routeExecute => routes_o(60), clock => clock, reset => reset);
	route_R62 : route_61 port map(routeRequest => routes_i(61), ne290_command => cmd_R62_ne290, track_ne290 => state_ne290, ne377_command => cmd_R62_ne377, track_ne377 => state_ne377, ne111_command => cmd_R62_ne111, track_ne111 => state_ne111, D14_command => cmd_R62_D14, D14_state => state_D14, D15_command => cmd_R62_D15, D15_state => state_D15, S86_state => state_S86, S86_command => cmd_R62_S86, T03_state => state_T03, T03_command =>cmd_R62_T03, routeExecute => routes_o(61), clock => clock, reset => reset);
	route_R63 : route_62 port map(routeRequest => routes_i(62), ne407_command => cmd_R63_ne407, track_ne407 => state_ne407, ne122_command => cmd_R63_ne122, track_ne122 => state_ne122, D16_command => cmd_R63_D16, D16_state => state_D16, S93_state => state_S93, S93_command => cmd_R63_S93, T17_state => state_T17, T17_command =>cmd_R63_T17, routeExecute => routes_o(62), clock => clock, reset => reset);
	route_R64 : route_63 port map(routeRequest => routes_i(63), ne61_command => cmd_R64_ne61, track_ne61 => state_ne61, ne407_command => cmd_R64_ne407, track_ne407 => state_ne407, ne98_command => cmd_R64_ne98, track_ne98 => state_ne98, ne99_command => cmd_R64_ne99, track_ne99 => state_ne99, ne123_command => cmd_R64_ne123, track_ne123 => state_ne123, Lc01_command => cmd_R64_Lc01, Lc01_state => state_Lc01, D08_command => cmd_R64_D08, D08_state => state_D08, D05_command => cmd_R64_D05, D05_state => state_D05, D16_command => cmd_R64_D16, D16_state => state_D16, S93_state => state_S93, S93_command => cmd_R64_S93, X51_state => state_X51, X51_command =>cmd_R64_X51, routeExecute => routes_o(63), clock => clock, reset => reset);
	route_R65 : route_64 port map(routeRequest => routes_i(64), ne63_command => cmd_R65_ne63, track_ne63 => state_ne63, ne65_command => cmd_R65_ne65, track_ne65 => state_ne65, D05_command => cmd_R65_D05, D05_state => state_D05, D18_command => cmd_R65_D18, D18_state => state_D18, C94_state => state_C94, C94_command => cmd_R65_C94, C54_state => state_C54, C54_command =>cmd_R65_C54, routeExecute => routes_o(64), clock => clock, reset => reset);
	route_R66 : route_65 port map(routeRequest => routes_i(65), ne63_command => cmd_R66_ne63, track_ne63 => state_ne63, ne65_command => cmd_R66_ne65, track_ne65 => state_ne65, D18_command => cmd_R66_D18, D18_state => state_D18, Sw01_command => cmd_R66_Sw01, Sw01_state => state_Sw01, S95_state => state_S95, S95_command => cmd_R66_S95, C119_state => state_C119, C119_command =>cmd_R66_C119, routeExecute => routes_o(65), clock => clock, reset => reset);
	route_R67 : route_66 port map(routeRequest => routes_i(66), ne63_command => cmd_R67_ne63, track_ne63 => state_ne63, ne421_command => cmd_R67_ne421, track_ne421 => state_ne421, ne124_command => cmd_R67_ne124, track_ne124 => state_ne124, D18_command => cmd_R67_D18, D18_state => state_D18, D19_command => cmd_R67_D19, D19_state => state_D19, S95_state => state_S95, S95_command => cmd_R67_S95, T05_state => state_T05, T05_command =>cmd_R67_T05, routeExecute => routes_o(66), clock => clock, reset => reset);
	route_R68 : route_67 port map(routeRequest => routes_i(67), ne114_command => cmd_R68_ne114, track_ne114 => state_ne114, ne132_command => cmd_R68_ne132, track_ne132 => state_ne132, D20_command => cmd_R68_D20, D20_state => state_D20, D23_command => cmd_R68_D23, D23_state => state_D23, S101_state => state_S101, S101_command => cmd_R68_S101, J47_state => state_J47, J47_command =>cmd_R68_J47, routeExecute => routes_o(67), clock => clock, reset => reset);
	route_R69 : route_68 port map(routeRequest => routes_i(68), ne114_command => cmd_R69_ne114, track_ne114 => state_ne114, ne127_command => cmd_R69_ne127, track_ne127 => state_ne127, ne129_command => cmd_R69_ne129, track_ne129 => state_ne129, D10_command => cmd_R69_D10, D10_state => state_D10, D09_command => cmd_R69_D09, D09_state => state_D09, D23_command => cmd_R69_D23, D23_state => state_D23, D24_command => cmd_R69_D24, D24_state => state_D24, D12_command => cmd_R69_D12, D12_state => state_D12, S101_state => state_S101, S101_command => cmd_R69_S101, S117_state => state_S117, S117_command =>cmd_R69_S117, routeExecute => routes_o(68), clock => clock, reset => reset);
	route_R70 : route_69 port map(routeRequest => routes_i(69), ne114_command => cmd_R70_ne114, track_ne114 => state_ne114, ne129_command => cmd_R70_ne129, track_ne129 => state_ne129, ne130_command => cmd_R70_ne130, track_ne130 => state_ne130, D10_command => cmd_R70_D10, D10_state => state_D10, D09_command => cmd_R70_D09, D09_state => state_D09, D23_command => cmd_R70_D23, D23_state => state_D23, D12_command => cmd_R70_D12, D12_state => state_D12, S101_state => state_S101, S101_command => cmd_R70_S101, C79_state => state_C79, C79_command =>cmd_R70_C79, routeExecute => routes_o(69), clock => clock, reset => reset);
	route_R71 : route_70 port map(routeRequest => routes_i(70), ne114_command => cmd_R71_ne114, track_ne114 => state_ne114, ne127_command => cmd_R71_ne127, track_ne127 => state_ne127, ne129_command => cmd_R71_ne129, track_ne129 => state_ne129, D23_command => cmd_R71_D23, D23_state => state_D23, D12_command => cmd_R71_D12, D12_state => state_D12, S104_state => state_S104, S104_command => cmd_R71_S104, L29_state => state_L29, L29_command =>cmd_R71_L29, routeExecute => routes_o(70), clock => clock, reset => reset);
	route_R72 : route_71 port map(routeRequest => routes_i(71), ne450_command => cmd_R72_ne450, track_ne450 => state_ne450, ne127_command => cmd_R72_ne127, track_ne127 => state_ne127, D12_command => cmd_R72_D12, D12_state => state_D12, S104_state => state_S104, S104_command => cmd_R72_S104, T07_state => state_T07, T07_command =>cmd_R72_T07, routeExecute => routes_o(71), clock => clock, reset => reset);
	route_R73 : route_72 port map(routeRequest => routes_i(72), ne114_command => cmd_R73_ne114, track_ne114 => state_ne114, ne129_command => cmd_R73_ne129, track_ne129 => state_ne129, ne130_command => cmd_R73_ne130, track_ne130 => state_ne130, D23_command => cmd_R73_D23, D23_state => state_D23, D12_command => cmd_R73_D12, D12_state => state_D12, S107_state => state_S107, S107_command => cmd_R73_S107, L29_state => state_L29, L29_command =>cmd_R73_L29, routeExecute => routes_o(72), clock => clock, reset => reset);
	route_R74 : route_73 port map(routeRequest => routes_i(73), ne450_command => cmd_R74_ne450, track_ne450 => state_ne450, ne130_command => cmd_R74_ne130, track_ne130 => state_ne130, D12_command => cmd_R74_D12, D12_state => state_D12, S107_state => state_S107, S107_command => cmd_R74_S107, T07_state => state_T07, T07_command =>cmd_R74_T07, routeExecute => routes_o(73), clock => clock, reset => reset);
	route_R75 : route_74 port map(routeRequest => routes_i(74), ne912_command => cmd_R75_ne912, track_ne912 => state_ne912, ne465_command => cmd_R75_ne465, track_ne465 => state_ne465, ne131_command => cmd_R75_ne131, track_ne131 => state_ne131, D20_command => cmd_R75_D20, D20_state => state_D20, D21_command => cmd_R75_D21, D21_state => state_D21, S110_state => state_S110, S110_command => cmd_R75_S110, T09_state => state_T09, T09_command =>cmd_R75_T09, routeExecute => routes_o(74), clock => clock, reset => reset);
	route_R76 : route_75 port map(routeRequest => routes_i(75), ne912_command => cmd_R76_ne912, track_ne912 => state_ne912, ne132_command => cmd_R76_ne132, track_ne132 => state_ne132, D20_command => cmd_R76_D20, D20_state => state_D20, D23_command => cmd_R76_D23, D23_state => state_D23, S110_state => state_S110, S110_command => cmd_R76_S110, J46_state => state_J46, J46_command =>cmd_R76_J46, routeExecute => routes_o(75), clock => clock, reset => reset);
	route_R77 : route_76 port map(routeRequest => routes_i(76), ne910_command => cmd_R77_ne910, track_ne910 => state_ne910, ne101_command => cmd_R77_ne101, track_ne101 => state_ne101, ne127_command => cmd_R77_ne127, track_ne127 => state_ne127, ne135_command => cmd_R77_ne135, track_ne135 => state_ne135, D10_command => cmd_R77_D10, D10_state => state_D10, D09_command => cmd_R77_D09, D09_state => state_D09, D24_command => cmd_R77_D24, D24_state => state_D24, S117_state => state_S117, S117_command => cmd_R77_S117, J43_state => state_J43, J43_command =>cmd_R77_J43, routeExecute => routes_o(76), clock => clock, reset => reset);
	route_R78 : route_77 port map(routeRequest => routes_i(77), ne127_command => cmd_R78_ne127, track_ne127 => state_ne127, ne134_command => cmd_R78_ne134, track_ne134 => state_ne134, D24_command => cmd_R78_D24, D24_state => state_D24, S117_state => state_S117, S117_command => cmd_R78_S117, T23_state => state_T23, T23_command =>cmd_R78_T23, routeExecute => routes_o(77), clock => clock, reset => reset);
	route_R79 : route_78 port map(routeRequest => routes_i(78), ne65_command => cmd_R79_ne65, track_ne65 => state_ne65, ne992_command => cmd_R79_ne992, track_ne992 => state_ne992, Sw01_command => cmd_R79_Sw01, Sw01_state => state_Sw01, C119_state => state_C119, C119_command => cmd_R79_C119, J40_state => state_J40, J40_command =>cmd_R79_J40, routeExecute => routes_o(78), clock => clock, reset => reset);
	route_R80 : route_79 port map(routeRequest => routes_i(79), ne65_command => cmd_R80_ne65, track_ne65 => state_ne65, ne992_command => cmd_R80_ne992, track_ne992 => state_ne992, D18_command => cmd_R80_D18, D18_state => state_D18, Sw01_command => cmd_R80_Sw01, Sw01_state => state_Sw01, S120_state => state_S120, S120_command => cmd_R80_S120, C94_state => state_C94, C94_command =>cmd_R80_C94, routeExecute => routes_o(79), clock => clock, reset => reset);
	route_R81 : route_80 port map(routeRequest => routes_i(80), ne400_command => cmd_R81_ne400, track_ne400 => state_ne400, ne992_command => cmd_R81_ne992, track_ne992 => state_ne992, ne994_command => cmd_R81_ne994, track_ne994 => state_ne994, Sw01_command => cmd_R81_Sw01, Sw01_state => state_Sw01, D07_command => cmd_R81_D07, D07_state => state_D07, Sw05_command => cmd_R81_Sw05, Sw05_state => state_Sw05, S120_state => state_S120, S120_command => cmd_R81_S120, S74_state => state_S74, S74_command =>cmd_R81_S74, routeExecute => routes_o(80), clock => clock, reset => reset);
	route_R82 : route_81 port map(routeRequest => routes_i(81), ne400_command => cmd_R82_ne400, track_ne400 => state_ne400, ne993_command => cmd_R82_ne993, track_ne993 => state_ne993, D07_command => cmd_R82_D07, D07_state => state_D07, Sw05_command => cmd_R82_Sw05, Sw05_state => state_Sw05, C122_state => state_C122, C122_command => cmd_R82_C122, S74_state => state_S74, S74_command =>cmd_R82_S74, routeExecute => routes_o(81), clock => clock, reset => reset);
	route_R83 : route_82 port map(routeRequest => routes_i(82), ne400_command => cmd_R83_ne400, track_ne400 => state_ne400, ne993_command => cmd_R83_ne993, track_ne993 => state_ne993, Sw05_command => cmd_R83_Sw05, Sw05_state => state_Sw05, S123_state => state_S123, S123_command => cmd_R83_S123, T25_state => state_T25, T25_command =>cmd_R83_T25, routeExecute => routes_o(82), clock => clock, reset => reset);
	route_R84 : route_83 port map(routeRequest => routes_i(83), ne400_command => cmd_R84_ne400, track_ne400 => state_ne400, ne992_command => cmd_R84_ne992, track_ne992 => state_ne992, ne994_command => cmd_R84_ne994, track_ne994 => state_ne994, Sw01_command => cmd_R84_Sw01, Sw01_state => state_Sw01, Sw05_command => cmd_R84_Sw05, Sw05_state => state_Sw05, S123_state => state_S123, S123_command => cmd_R84_S123, J40_state => state_J40, J40_command =>cmd_R84_J40, routeExecute => routes_o(83), clock => clock, reset => reset);
	route_R85 : route_84 port map(routeRequest => routes_i(84), ne297_command => cmd_R85_ne297, track_ne297 => state_ne297, ne995_command => cmd_R85_ne995, track_ne995 => state_ne995, D04_command => cmd_R85_D04, D04_state => state_D04, Sw03_command => cmd_R85_Sw03, Sw03_state => state_Sw03, C125_state => state_C125, C125_command => cmd_R85_C125, S71_state => state_S71, S71_command =>cmd_R85_S71, routeExecute => routes_o(84), clock => clock, reset => reset);
	route_R86 : route_85 port map(routeRequest => routes_i(85), ne297_command => cmd_R86_ne297, track_ne297 => state_ne297, ne995_command => cmd_R86_ne995, track_ne995 => state_ne995, Sw03_command => cmd_R86_Sw03, Sw03_state => state_Sw03, S126_state => state_S126, S126_command => cmd_R86_S126, T27_state => state_T27, T27_command =>cmd_R86_T27, routeExecute => routes_o(85), clock => clock, reset => reset);
	route_R87 : route_86 port map(routeRequest => routes_i(86), ne297_command => cmd_R87_ne297, track_ne297 => state_ne297, ne996_command => cmd_R87_ne996, track_ne996 => state_ne996, ne997_command => cmd_R87_ne997, track_ne997 => state_ne997, Sw04_command => cmd_R87_Sw04, Sw04_state => state_Sw04, Sw03_command => cmd_R87_Sw03, Sw03_state => state_Sw03, S126_state => state_S126, S126_command => cmd_R87_S126, J38_state => state_J38, J38_command =>cmd_R87_J38, routeExecute => routes_o(86), clock => clock, reset => reset);
	route_R88 : route_87 port map(routeRequest => routes_i(87), ne292_command => cmd_R88_ne292, track_ne292 => state_ne292, ne996_command => cmd_R88_ne996, track_ne996 => state_ne996, D14_command => cmd_R88_D14, D14_state => state_D14, Sw04_command => cmd_R88_Sw04, Sw04_state => state_Sw04, S129_state => state_S129, S129_command => cmd_R88_S129, J37_state => state_J37, J37_command =>cmd_R88_J37, routeExecute => routes_o(87), clock => clock, reset => reset);
	route_R89 : route_88 port map(routeRequest => routes_i(88), ne297_command => cmd_R89_ne297, track_ne297 => state_ne297, ne996_command => cmd_R89_ne996, track_ne996 => state_ne996, ne997_command => cmd_R89_ne997, track_ne997 => state_ne997, Sw04_command => cmd_R89_Sw04, Sw04_state => state_Sw04, D04_command => cmd_R89_D04, D04_state => state_D04, Sw03_command => cmd_R89_Sw03, Sw03_state => state_Sw03, S129_state => state_S129, S129_command => cmd_R89_S129, S71_state => state_S71, S71_command =>cmd_R89_S71, routeExecute => routes_o(88), clock => clock, reset => reset);
	processed <= processing;
	tracks_o(0) <= state_ne991;
	tracks_o(1) <= state_ne61;
	tracks_o(2) <= state_ne63;
	tracks_o(3) <= state_ne65;
	tracks_o(4) <= state_ne910;
	tracks_o(5) <= state_ne912;
	tracks_o(6) <= state_ne114;
	tracks_o(7) <= state_ne288;
	tracks_o(8) <= state_ne290;
	tracks_o(9) <= state_ne292;
	tracks_o(10) <= state_ne295;
	tracks_o(11) <= state_ne297;
	tracks_o(12) <= state_ne377;
	tracks_o(13) <= state_ne384;
	tracks_o(14) <= state_ne400;
	tracks_o(15) <= state_ne404;
	tracks_o(16) <= state_ne407;
	tracks_o(17) <= state_ne421;
	tracks_o(18) <= state_ne450;
	tracks_o(19) <= state_ne465;
	tracks_o(20) <= state_ne98;
	tracks_o(21) <= state_ne99;
	tracks_o(22) <= state_ne100;
	tracks_o(23) <= state_ne101;
	tracks_o(24) <= state_ne102;
	tracks_o(25) <= state_ne104;
	tracks_o(26) <= state_ne110;
	tracks_o(27) <= state_ne111;
	tracks_o(28) <= state_ne113;
	tracks_o(29) <= state_ne122;
	tracks_o(30) <= state_ne123;
	tracks_o(31) <= state_ne124;
	tracks_o(32) <= state_ne126;
	tracks_o(33) <= state_ne127;
	tracks_o(34) <= state_ne129;
	tracks_o(35) <= state_ne130;
	tracks_o(36) <= state_ne131;
	tracks_o(37) <= state_ne132;
	tracks_o(38) <= state_ne133;
	tracks_o(39) <= state_ne134;
	tracks_o(40) <= state_ne135;
	tracks_o(41) <= state_ne992;
	tracks_o(42) <= state_ne993;
	tracks_o(43) <= state_ne994;
	tracks_o(44) <= state_ne995;
	tracks_o(45) <= state_ne996;
	tracks_o(46) <= state_ne997;
end Behavioral;