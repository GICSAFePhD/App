--  route_48.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity route_48 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne384_state : in nodeStates;
			ne384_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_command : out routeCommands;
			ne288_state : in nodeStates;
			ne288_command : out routeCommands;
			ne991_state : in nodeStates;
			ne991_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_command : out routeCommands;
			routeState : out std_logic
		);
	end entity route_48;
architecture Behavioral of route_48 is
begin
	routeState <= '0';
end Behavioral;