--  network.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity network is
		generic(
			N : natural := 316;
			N_SIGNALS : natural := 77;
			N_ROUTES : natural := 89;
			N_LEVELCROSSINGS : natural := 2;
			N_SINGLESWITCHES : natural := 22;
			N_DOUBLEWITCHES : natural := 1;
			N_TRACKCIRCUITS : natural := 47
		);
		port(
			clock : in std_logic;
			processing : in std_logic;
			processed : out std_logic;
			ocupation : in std_logic_vector(N_TRACKCIRCUITS-1 downto 0);
			signals_i : in signals_type;
			signals_o : out signals_type;
			routes_i : in std_logic_vector(N_ROUTES-1 downto 0);
			routes_o : out std_logic_vector(N_ROUTES-1 downto 0);
			levelCrossings_i : in std_logic_vector(N_LEVELCROSSINGS-1 downto 0);
			levelCrossings_o : out std_logic_vector(N_LEVELCROSSINGS-1 downto 0);
			singleSwitches_i : in std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			singleSwitches_o : out std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			doubleSwitches_i : in dSwitch_type;
			doubleSwitches_o : out dSwitch_type;
			reset : in std_logic
		);
	end entity network;
architecture Behavioral of network is
	component levelCrossing_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation_ne98 : in std_logic;
			ocupation_ne996 : in std_logic;
			ocupation_ne99 : in std_logic;
			R30_command : in routeCommands;
			R31_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc01 : out levelCrossingStates;
			lock_Lc01 : out objectLock
		);
	end component levelCrossing_0;
	component levelCrossing_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne992 : in std_logic;
			ocupation_ne101 : in std_logic;
			R32_command : in routeCommands;
			R33_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc04 : out levelCrossingStates;
			lock_Lc04 : out objectLock
		);
	end component levelCrossing_1;
	component singleSwitch_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R20_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			R41_command : in routeCommands;
			R60_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D01 : out singleSwitchStates;
			lock_D01 : out objectLock
		);
	end component singleSwitch_0;
	component singleSwitch_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R51_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R64_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D08 : out singleSwitchStates;
			lock_D08 : out objectLock
		);
	end component singleSwitch_1;
	component singleSwitch_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R34_command : in routeCommands;
			R35_command : in routeCommands;
			R36_command : in routeCommands;
			R51_command : in routeCommands;
			R64_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D05 : out singleSwitchStates;
			lock_D05 : out objectLock
		);
	end component singleSwitch_2;
	component singleSwitch_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R67_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D18 : out singleSwitchStates;
			lock_D18 : out objectLock
		);
	end component singleSwitch_3;
	component singleSwitch_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			R81_command : in routeCommands;
			R84_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw01 : out singleSwitchStates;
			lock_Sw01 : out objectLock
		);
	end component singleSwitch_4;
	component singleSwitch_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			R58_command : in routeCommands;
			R77_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D10 : out singleSwitchStates;
			lock_D10 : out objectLock
		);
	end component singleSwitch_5;
	component singleSwitch_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R26_command : in routeCommands;
			R37_command : in routeCommands;
			R38_command : in routeCommands;
			R55_command : in routeCommands;
			R77_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D09 : out singleSwitchStates;
			lock_D09 : out objectLock
		);
	end component singleSwitch_6;
	component singleSwitch_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R8_command : in routeCommands;
			R28_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D20 : out singleSwitchStates;
			lock_D20 : out objectLock
		);
	end component singleSwitch_7;
	component singleSwitch_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R27_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R73_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D23 : out singleSwitchStates;
			lock_D23 : out objectLock
		);
	end component singleSwitch_8;
	component singleSwitch_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			R60_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D03 : out singleSwitchStates;
			lock_D03 : out objectLock
		);
	end component singleSwitch_9;
	component singleSwitch_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R2_command : in routeCommands;
			R22_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D14 : out singleSwitchStates;
			lock_D14 : out objectLock
		);
	end component singleSwitch_10;
	component singleSwitch_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R21_command : in routeCommands;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			R89_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw04 : out singleSwitchStates;
			lock_Sw04 : out objectLock
		);
	end component singleSwitch_11;
	component singleSwitch_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R11_command : in routeCommands;
			R42_command : in routeCommands;
			R45_command : in routeCommands;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D04 : out singleSwitchStates;
			lock_D04 : out objectLock
		);
	end component singleSwitch_12;
	component singleSwitch_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			R87_command : in routeCommands;
			R89_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw03 : out singleSwitchStates;
			lock_Sw03 : out objectLock
		);
	end component singleSwitch_13;
	component singleSwitch_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R2_command : in routeCommands;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			R62_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D15 : out singleSwitchStates;
			lock_D15 : out objectLock
		);
	end component singleSwitch_14;
	component singleSwitch_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R11_command : in routeCommands;
			R42_command : in routeCommands;
			R59_command : in routeCommands;
			R60_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw02 : out singleSwitchStates;
			lock_Sw02 : out objectLock
		);
	end component singleSwitch_15;
	component singleSwitch_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R13_command : in routeCommands;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			R52_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D07 : out singleSwitchStates;
			lock_D07 : out objectLock
		);
	end component singleSwitch_16;
	component singleSwitch_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R81_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			R84_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw05 : out singleSwitchStates;
			lock_Sw05 : out objectLock
		);
	end component singleSwitch_17;
	component singleSwitch_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R13_command : in routeCommands;
			R52_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D16 : out singleSwitchStates;
			lock_D16 : out objectLock
		);
	end component singleSwitch_18;
	component singleSwitch_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			R67_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D19 : out singleSwitchStates;
			lock_D19 : out objectLock
		);
	end component singleSwitch_19;
	component singleSwitch_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R8_command : in routeCommands;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			R75_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D21 : out singleSwitchStates;
			lock_D21 : out objectLock
		);
	end component singleSwitch_20;
	component singleSwitch_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R16_command : in routeCommands;
			R56_command : in routeCommands;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_D24 : out singleSwitchStates;
			lock_D24 : out objectLock
		);
	end component singleSwitch_21;
	component doubleSwitch_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R6_command : in routeCommands;
			R7_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			indication : in dSwitch_type;
			command : out dSwitch_type;
			correspondence_D12 : out doubleSwitchStates;
			lock_D12 : out objectLock
		);
	end component doubleSwitch_0;
	component railwaySignal_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne991 : in std_logic;
			correspondence_T01 : out signalStates;
			lock_T01 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_0;
	component railwaySignal_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R1_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne991 : in std_logic;
			correspondence_T02 : out signalStates;
			lock_T02 : out objectLock;
			correspondence_S64 : in signalStates;
			--Ocupation level 2
			ocupation_ne290 : in std_logic;
			ocupation_ne288 : in std_logic;
			correspondence_S69 : in signalStates;
			correspondence_S86 : in signalStates;
			D01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_1;
	component railwaySignal_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne991 : in std_logic;
			correspondence_S64 : out signalStates;
			lock_S64 : out objectLock;
			--Ocupation level 1
			ocupation_ne288 : in std_logic;
			ocupation_ne290 : in std_logic;
			correspondence_S69 : in signalStates;
			correspondence_S86 : in signalStates;
			D01_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne110 : in std_logic;
			ocupation_ne295 : in std_logic;
			ocupation_ne111 : in std_logic;
			ocupation_ne377 : in std_logic;
			ocupation_ne292 : in std_logic;
			correspondence_C70 : in signalStates;
			correspondence_B68 : in signalStates;
			correspondence_J36 : in signalStates;
			correspondence_T03 : in signalStates;
			D03_state : in singleSwitchStates;
			D14_state : in singleSwitchStates;
			D15_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_2;
	component railwaySignal_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne61 : in std_logic;
			correspondence_S78 : out signalStates;
			lock_S78 : out objectLock;
			--Ocupation level 1
			ocupation_ne404 : in std_logic;
			ocupation_ne123 : in std_logic;
			correspondence_C73 : in signalStates;
			correspondence_B77 : in signalStates;
			D08_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne400 : in std_logic;
			ocupation_ne407 : in std_logic;
			correspondence_S123 : in signalStates;
			D07_state : in singleSwitchStates;
			D16_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_3;
	component railwaySignal_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R34_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne63 : in std_logic;
			correspondence_C54 : out signalStates;
			lock_C54 : out objectLock;
			--Ocupation level 1
			ocupation_ne99 : in std_logic;
			ocupation_ne98 : in std_logic;
			correspondence_X51 : in signalStates;
			D05_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne996 : in std_logic;
			correspondence_S129 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_4;
	component railwaySignal_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R66_command : in routeCommands;
			R67_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne63 : in std_logic;
			correspondence_S95 : out signalStates;
			lock_S95 : out objectLock;
			--Ocupation level 1
			ocupation_ne65 : in std_logic;
			ocupation_ne124 : in std_logic;
			ocupation_ne421 : in std_logic;
			correspondence_C119 : in signalStates;
			correspondence_T05 : in signalStates;
			D18_state : in singleSwitchStates;
			D19_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne992 : in std_logic;
			correspondence_J40 : in signalStates;
			Sw01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_5;
	component railwaySignal_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R65_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne65 : in std_logic;
			correspondence_C94 : out signalStates;
			lock_C94 : out objectLock;
			--Ocupation level 1
			ocupation_ne63 : in std_logic;
			correspondence_C54 : in signalStates;
			D18_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne98 : in std_logic;
			ocupation_ne99 : in std_logic;
			correspondence_X51 : in signalStates;
			D05_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_6;
	component railwaySignal_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R79_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne65 : in std_logic;
			correspondence_C119 : out signalStates;
			lock_C119 : out objectLock;
			--Ocupation level 1
			ocupation_ne992 : in std_logic;
			correspondence_J40 : in signalStates;
			Sw01_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne100 : in std_logic;
			correspondence_L31 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_7;
	component railwaySignal_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R57_command : in routeCommands;
			R58_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne910 : in std_logic;
			correspondence_S81 : out signalStates;
			lock_S81 : out objectLock;
			--Ocupation level 1
			ocupation_ne130 : in std_logic;
			ocupation_ne135 : in std_logic;
			correspondence_S107 : in signalStates;
			correspondence_B80 : in signalStates;
			D10_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne114 : in std_logic;
			ocupation_ne450 : in std_logic;
			ocupation_ne129 : in std_logic;
			ocupation_ne127 : in std_logic;
			correspondence_L29 : in signalStates;
			correspondence_T07 : in signalStates;
			correspondence_S104 : in signalStates;
			D23_state : in singleSwitchStates;
			D12_state : in doubleSwitchStates;
			D24_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_8;
	component railwaySignal_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R26_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne912 : in std_logic;
			correspondence_J45 : out signalStates;
			lock_J45 : out objectLock;
			--Ocupation level 1
			ocupation_ne101 : in std_logic;
			correspondence_J43 : in signalStates;
			D09_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne100 : in std_logic;
			correspondence_X53 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_9;
	component railwaySignal_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne912 : in std_logic;
			correspondence_S110 : out signalStates;
			lock_S110 : out objectLock;
			--Ocupation level 1
			ocupation_ne131 : in std_logic;
			ocupation_ne465 : in std_logic;
			ocupation_ne132 : in std_logic;
			correspondence_T09 : in signalStates;
			correspondence_J46 : in signalStates;
			D20_state : in singleSwitchStates;
			D21_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne114 : in std_logic;
			correspondence_L29 : in signalStates;
			D23_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_10;
	component railwaySignal_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R17_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne114 : in std_logic;
			correspondence_L29 : out signalStates;
			lock_L29 : out objectLock;
			correspondence_J48 : in signalStates;
			--Ocupation level 2
			ocupation_ne102 : in std_logic;
			correspondence_T11 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_11;
	component railwaySignal_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R29_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne114 : in std_logic;
			correspondence_J48 : out signalStates;
			lock_J48 : out objectLock;
			--Ocupation level 1
			ocupation_ne102 : in std_logic;
			correspondence_T11 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_12;
	component railwaySignal_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne114 : in std_logic;
			correspondence_S101 : out signalStates;
			lock_S101 : out objectLock;
			--Ocupation level 1
			ocupation_ne132 : in std_logic;
			ocupation_ne129 : in std_logic;
			ocupation_ne127 : in std_logic;
			ocupation_ne130 : in std_logic;
			correspondence_J47 : in signalStates;
			correspondence_S117 : in signalStates;
			correspondence_C79 : in signalStates;
			D23_state : in singleSwitchStates;
			D12_state : in doubleSwitchStates;
			--Ocupation level 2
			ocupation_ne912 : in std_logic;
			ocupation_ne910 : in std_logic;
			ocupation_ne134 : in std_logic;
			ocupation_ne135 : in std_logic;
			ocupation_ne101 : in std_logic;
			correspondence_J45 : in signalStates;
			correspondence_J43 : in signalStates;
			correspondence_T23 : in signalStates;
			D20_state : in singleSwitchStates;
			D09_state : in singleSwitchStates;
			D10_state : in singleSwitchStates;
			D24_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_13;
	component railwaySignal_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne288 : in std_logic;
			correspondence_S69 : out signalStates;
			lock_S69 : out objectLock;
			--Ocupation level 1
			ocupation_ne295 : in std_logic;
			ocupation_ne110 : in std_logic;
			correspondence_C70 : in signalStates;
			correspondence_B68 : in signalStates;
			D03_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne297 : in std_logic;
			ocupation_ne384 : in std_logic;
			correspondence_S126 : in signalStates;
			D04_state : in singleSwitchStates;
			Sw02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_14;
	component railwaySignal_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R20_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne290 : in std_logic;
			correspondence_J35 : out signalStates;
			lock_J35 : out objectLock;
			--Ocupation level 1
			ocupation_ne991 : in std_logic;
			correspondence_T01 : in signalStates;
			D01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_15;
	component railwaySignal_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne290 : in std_logic;
			correspondence_S86 : out signalStates;
			lock_S86 : out objectLock;
			--Ocupation level 1
			ocupation_ne292 : in std_logic;
			ocupation_ne111 : in std_logic;
			ocupation_ne377 : in std_logic;
			correspondence_J36 : in signalStates;
			correspondence_T03 : in signalStates;
			D14_state : in singleSwitchStates;
			D15_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne996 : in std_logic;
			correspondence_J38 : in signalStates;
			Sw04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_16;
	component railwaySignal_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R21_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne292 : in std_logic;
			correspondence_J36 : out signalStates;
			lock_J36 : out objectLock;
			--Ocupation level 1
			ocupation_ne996 : in std_logic;
			correspondence_J38 : in signalStates;
			Sw04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne98 : in std_logic;
			correspondence_L30 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_17;
	component railwaySignal_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R22_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne292 : in std_logic;
			correspondence_J37 : out signalStates;
			lock_J37 : out objectLock;
			--Ocupation level 1
			ocupation_ne290 : in std_logic;
			correspondence_J35 : in signalStates;
			D14_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne991 : in std_logic;
			correspondence_T01 : in signalStates;
			D01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_18;
	component railwaySignal_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R41_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne295 : in std_logic;
			correspondence_C67 : out signalStates;
			lock_C67 : out objectLock;
			--Ocupation level 1
			ocupation_ne288 : in std_logic;
			ocupation_ne991 : in std_logic;
			correspondence_T01 : in signalStates;
			D01_state : in singleSwitchStates;
			D03_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_19;
	component railwaySignal_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R45_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne295 : in std_logic;
			correspondence_C70 : out signalStates;
			lock_C70 : out objectLock;
			--Ocupation level 1
			ocupation_ne297 : in std_logic;
			correspondence_S126 : in signalStates;
			D04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne996 : in std_logic;
			ocupation_ne995 : in std_logic;
			ocupation_ne997 : in std_logic;
			correspondence_T27 : in signalStates;
			correspondence_J38 : in signalStates;
			Sw03_state : in singleSwitchStates;
			Sw04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_20;
	component railwaySignal_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne297 : in std_logic;
			correspondence_S71 : out signalStates;
			lock_S71 : out objectLock;
			--Ocupation level 1
			ocupation_ne295 : in std_logic;
			ocupation_ne384 : in std_logic;
			correspondence_C67 : in signalStates;
			correspondence_S84 : in signalStates;
			D04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne991 : in std_logic;
			ocupation_ne288 : in std_logic;
			ocupation_ne110 : in std_logic;
			ocupation_ne104 : in std_logic;
			correspondence_T01 : in signalStates;
			correspondence_T13 : in signalStates;
			D01_state : in singleSwitchStates;
			D03_state : in singleSwitchStates;
			Sw02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_21;
	component railwaySignal_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R86_command : in routeCommands;
			R87_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne297 : in std_logic;
			correspondence_S126 : out signalStates;
			lock_S126 : out objectLock;
			--Ocupation level 1
			ocupation_ne995 : in std_logic;
			ocupation_ne997 : in std_logic;
			ocupation_ne996 : in std_logic;
			correspondence_T27 : in signalStates;
			correspondence_J38 : in signalStates;
			Sw03_state : in singleSwitchStates;
			Sw04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne98 : in std_logic;
			correspondence_L30 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_22;
	component railwaySignal_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne377 : in std_logic;
			correspondence_T03 : out signalStates;
			lock_T03 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_23;
	component railwaySignal_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R2_command : in routeCommands;
			R3_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne377 : in std_logic;
			correspondence_T04 : out signalStates;
			lock_T04 : out objectLock;
			--Ocupation level 1
			ocupation_ne111 : in std_logic;
			ocupation_ne290 : in std_logic;
			ocupation_ne113 : in std_logic;
			correspondence_J35 : in signalStates;
			correspondence_T15 : in signalStates;
			D14_state : in singleSwitchStates;
			D15_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne991 : in std_logic;
			correspondence_T01 : in signalStates;
			D01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_24;
	component railwaySignal_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R59_command : in routeCommands;
			R60_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne384 : in std_logic;
			correspondence_S84 : out signalStates;
			lock_S84 : out objectLock;
			--Ocupation level 1
			ocupation_ne104 : in std_logic;
			ocupation_ne110 : in std_logic;
			ocupation_ne288 : in std_logic;
			ocupation_ne991 : in std_logic;
			correspondence_T13 : in signalStates;
			correspondence_T01 : in signalStates;
			Sw02_state : in singleSwitchStates;
			D01_state : in singleSwitchStates;
			D03_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_25;
	component railwaySignal_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne400 : in std_logic;
			correspondence_S74 : out signalStates;
			lock_S74 : out objectLock;
			--Ocupation level 1
			ocupation_ne404 : in std_logic;
			ocupation_ne407 : in std_logic;
			correspondence_C76 : in signalStates;
			correspondence_S93 : in signalStates;
			D07_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne98 : in std_logic;
			ocupation_ne99 : in std_logic;
			ocupation_ne61 : in std_logic;
			ocupation_ne123 : in std_logic;
			ocupation_ne122 : in std_logic;
			correspondence_X51 : in signalStates;
			correspondence_T17 : in signalStates;
			D05_state : in singleSwitchStates;
			D08_state : in singleSwitchStates;
			D16_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_26;
	component railwaySignal_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R83_command : in routeCommands;
			R84_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne400 : in std_logic;
			correspondence_S123 : out signalStates;
			lock_S123 : out objectLock;
			--Ocupation level 1
			ocupation_ne993 : in std_logic;
			ocupation_ne994 : in std_logic;
			ocupation_ne992 : in std_logic;
			correspondence_T25 : in signalStates;
			correspondence_J40 : in signalStates;
			Sw05_state : in singleSwitchStates;
			Sw01_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne100 : in std_logic;
			correspondence_L31 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_27;
	component railwaySignal_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R48_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne404 : in std_logic;
			correspondence_C73 : out signalStates;
			lock_C73 : out objectLock;
			--Ocupation level 1
			ocupation_ne400 : in std_logic;
			correspondence_S123 : in signalStates;
			D07_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne992 : in std_logic;
			ocupation_ne994 : in std_logic;
			ocupation_ne993 : in std_logic;
			correspondence_T25 : in signalStates;
			correspondence_J40 : in signalStates;
			Sw05_state : in singleSwitchStates;
			Sw01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_28;
	component railwaySignal_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R51_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne404 : in std_logic;
			correspondence_C76 : out signalStates;
			lock_C76 : out objectLock;
			--Ocupation level 1
			ocupation_ne61 : in std_logic;
			ocupation_ne99 : in std_logic;
			ocupation_ne98 : in std_logic;
			correspondence_X51 : in signalStates;
			D05_state : in singleSwitchStates;
			D08_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne996 : in std_logic;
			correspondence_S129 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_29;
	component railwaySignal_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne407 : in std_logic;
			correspondence_S93 : out signalStates;
			lock_S93 : out objectLock;
			--Ocupation level 1
			ocupation_ne122 : in std_logic;
			ocupation_ne123 : in std_logic;
			ocupation_ne61 : in std_logic;
			ocupation_ne99 : in std_logic;
			ocupation_ne98 : in std_logic;
			correspondence_T17 : in signalStates;
			correspondence_X51 : in signalStates;
			D16_state : in singleSwitchStates;
			D05_state : in singleSwitchStates;
			D08_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne996 : in std_logic;
			correspondence_S129 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_30;
	component railwaySignal_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne421 : in std_logic;
			correspondence_T05 : out signalStates;
			lock_T05 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_31;
	component railwaySignal_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			R5_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne421 : in std_logic;
			correspondence_T06 : out signalStates;
			lock_T06 : out objectLock;
			--Ocupation level 1
			ocupation_ne124 : in std_logic;
			ocupation_ne63 : in std_logic;
			ocupation_ne126 : in std_logic;
			correspondence_C54 : in signalStates;
			correspondence_T19 : in signalStates;
			D18_state : in singleSwitchStates;
			D19_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne98 : in std_logic;
			ocupation_ne99 : in std_logic;
			correspondence_X51 : in signalStates;
			D05_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_32;
	component railwaySignal_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne450 : in std_logic;
			correspondence_T07 : out signalStates;
			lock_T07 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_33;
	component railwaySignal_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R6_command : in routeCommands;
			R7_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne450 : in std_logic;
			correspondence_T08 : out signalStates;
			lock_T08 : out objectLock;
			--Ocupation level 1
			ocupation_ne127 : in std_logic;
			ocupation_ne130 : in std_logic;
			correspondence_S117 : in signalStates;
			correspondence_C79 : in signalStates;
			D12_state : in doubleSwitchStates;
			--Ocupation level 2
			ocupation_ne910 : in std_logic;
			ocupation_ne134 : in std_logic;
			ocupation_ne135 : in std_logic;
			ocupation_ne101 : in std_logic;
			correspondence_J43 : in signalStates;
			correspondence_T23 : in signalStates;
			D09_state : in singleSwitchStates;
			D10_state : in singleSwitchStates;
			D24_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_34;
	component railwaySignal_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne465 : in std_logic;
			correspondence_T09 : out signalStates;
			lock_T09 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_35;
	component railwaySignal_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R8_command : in routeCommands;
			R9_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne465 : in std_logic;
			correspondence_T10 : out signalStates;
			lock_T10 : out objectLock;
			--Ocupation level 1
			ocupation_ne131 : in std_logic;
			ocupation_ne912 : in std_logic;
			ocupation_ne133 : in std_logic;
			correspondence_J45 : in signalStates;
			correspondence_T21 : in signalStates;
			D20_state : in singleSwitchStates;
			D21_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne101 : in std_logic;
			correspondence_J43 : in signalStates;
			D09_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_36;
	component railwaySignal_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R18_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne98 : in std_logic;
			correspondence_L30 : out signalStates;
			lock_L30 : out objectLock;
			correspondence_X50 : in signalStates;
			--Ocupation level 2
			ocupation_ne99 : in std_logic;
			correspondence_S55 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_37;
	component railwaySignal_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R30_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne98 : in std_logic;
			correspondence_X50 : out signalStates;
			lock_X50 : out objectLock;
			--Ocupation level 1
			ocupation_ne99 : in std_logic;
			correspondence_S55 : in signalStates;
			--Ocupation level 2
			ocupation_ne61 : in std_logic;
			ocupation_ne63 : in std_logic;
			correspondence_S78 : in signalStates;
			correspondence_S95 : in signalStates;
			D05_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_38;
	component railwaySignal_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R31_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne98 : in std_logic;
			correspondence_X51 : out signalStates;
			lock_X51 : out objectLock;
			--Ocupation level 1
			ocupation_ne996 : in std_logic;
			correspondence_S129 : in signalStates;
			--Ocupation level 2
			ocupation_ne297 : in std_logic;
			ocupation_ne292 : in std_logic;
			ocupation_ne997 : in std_logic;
			correspondence_J37 : in signalStates;
			correspondence_S71 : in signalStates;
			Sw04_state : in singleSwitchStates;
			Sw03_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_39;
	component railwaySignal_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R35_command : in routeCommands;
			R36_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne99 : in std_logic;
			correspondence_S55 : out signalStates;
			lock_S55 : out objectLock;
			--Ocupation level 1
			ocupation_ne61 : in std_logic;
			ocupation_ne63 : in std_logic;
			correspondence_S78 : in signalStates;
			correspondence_S95 : in signalStates;
			D05_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne123 : in std_logic;
			ocupation_ne404 : in std_logic;
			ocupation_ne421 : in std_logic;
			ocupation_ne65 : in std_logic;
			ocupation_ne124 : in std_logic;
			correspondence_C73 : in signalStates;
			correspondence_B77 : in signalStates;
			correspondence_C119 : in signalStates;
			correspondence_T05 : in signalStates;
			D08_state : in singleSwitchStates;
			D18_state : in singleSwitchStates;
			D19_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_40;
	component railwaySignal_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R19_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne100 : in std_logic;
			correspondence_L31 : out signalStates;
			lock_L31 : out objectLock;
			correspondence_X52 : in signalStates;
			--Ocupation level 2
			ocupation_ne101 : in std_logic;
			correspondence_S59 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_41;
	component railwaySignal_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R32_command : in routeCommands;
			Lc04_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne100 : in std_logic;
			correspondence_X52 : out signalStates;
			lock_X52 : out objectLock;
			--Ocupation level 1
			ocupation_ne101 : in std_logic;
			correspondence_S59 : in signalStates;
			--Ocupation level 2
			ocupation_ne910 : in std_logic;
			ocupation_ne912 : in std_logic;
			correspondence_S110 : in signalStates;
			correspondence_S81 : in signalStates;
			D09_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_42;
	component railwaySignal_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R33_command : in routeCommands;
			Lc04_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne100 : in std_logic;
			correspondence_X53 : out signalStates;
			lock_X53 : out objectLock;
			--Ocupation level 1
			ocupation_ne992 : in std_logic;
			correspondence_S120 : in signalStates;
			--Ocupation level 2
			ocupation_ne65 : in std_logic;
			ocupation_ne994 : in std_logic;
			ocupation_ne400 : in std_logic;
			correspondence_C94 : in signalStates;
			correspondence_S74 : in signalStates;
			Sw01_state : in singleSwitchStates;
			Sw05_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_43;
	component railwaySignal_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R25_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne101 : in std_logic;
			correspondence_J43 : out signalStates;
			lock_J43 : out objectLock;
			--Ocupation level 1
			ocupation_ne100 : in std_logic;
			correspondence_X53 : in signalStates;
			--Ocupation level 2
			ocupation_ne992 : in std_logic;
			correspondence_S120 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_44;
	component railwaySignal_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R37_command : in routeCommands;
			R38_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne101 : in std_logic;
			correspondence_S59 : out signalStates;
			lock_S59 : out objectLock;
			--Ocupation level 1
			ocupation_ne912 : in std_logic;
			ocupation_ne910 : in std_logic;
			correspondence_S110 : in signalStates;
			correspondence_S81 : in signalStates;
			D09_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne132 : in std_logic;
			ocupation_ne465 : in std_logic;
			ocupation_ne131 : in std_logic;
			ocupation_ne130 : in std_logic;
			ocupation_ne135 : in std_logic;
			correspondence_T09 : in signalStates;
			correspondence_J46 : in signalStates;
			correspondence_S107 : in signalStates;
			correspondence_B80 : in signalStates;
			D20_state : in singleSwitchStates;
			D21_state : in singleSwitchStates;
			D10_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_45;
	component railwaySignal_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne102 : in std_logic;
			correspondence_T11 : out signalStates;
			lock_T11 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_46;
	component railwaySignal_47 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R10_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne102 : in std_logic;
			correspondence_T12 : out signalStates;
			lock_T12 : out objectLock;
			--Ocupation level 1
			ocupation_ne114 : in std_logic;
			correspondence_S101 : in signalStates;
			--Ocupation level 2
			ocupation_ne132 : in std_logic;
			ocupation_ne130 : in std_logic;
			ocupation_ne127 : in std_logic;
			ocupation_ne129 : in std_logic;
			correspondence_J47 : in signalStates;
			correspondence_S117 : in signalStates;
			correspondence_C79 : in signalStates;
			D23_state : in singleSwitchStates;
			D12_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_47;
	component railwaySignal_48 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne104 : in std_logic;
			correspondence_T13 : out signalStates;
			lock_T13 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_48;
	component railwaySignal_49 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R11_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne104 : in std_logic;
			correspondence_T14 : out signalStates;
			lock_T14 : out objectLock;
			--Ocupation level 1
			ocupation_ne384 : in std_logic;
			ocupation_ne297 : in std_logic;
			correspondence_S126 : in signalStates;
			D04_state : in singleSwitchStates;
			Sw02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne996 : in std_logic;
			ocupation_ne995 : in std_logic;
			ocupation_ne997 : in std_logic;
			correspondence_T27 : in signalStates;
			correspondence_J38 : in signalStates;
			Sw03_state : in singleSwitchStates;
			Sw04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_49;
	component railwaySignal_50 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R42_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne110 : in std_logic;
			correspondence_B68 : out signalStates;
			lock_B68 : out objectLock;
			--Ocupation level 1
			ocupation_ne384 : in std_logic;
			ocupation_ne297 : in std_logic;
			correspondence_S126 : in signalStates;
			D04_state : in singleSwitchStates;
			Sw02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne996 : in std_logic;
			ocupation_ne995 : in std_logic;
			ocupation_ne997 : in std_logic;
			correspondence_T27 : in signalStates;
			correspondence_J38 : in signalStates;
			Sw03_state : in singleSwitchStates;
			Sw04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_50;
	component railwaySignal_51 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne113 : in std_logic;
			correspondence_T15 : out signalStates;
			lock_T15 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_51;
	component railwaySignal_52 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R12_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne113 : in std_logic;
			correspondence_T16 : out signalStates;
			lock_T16 : out objectLock;
			--Ocupation level 1
			ocupation_ne377 : in std_logic;
			correspondence_T03 : in signalStates;
			D15_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_52;
	component railwaySignal_53 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne122 : in std_logic;
			correspondence_T17 : out signalStates;
			lock_T17 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_53;
	component railwaySignal_54 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R13_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne122 : in std_logic;
			correspondence_T18 : out signalStates;
			lock_T18 : out objectLock;
			--Ocupation level 1
			ocupation_ne407 : in std_logic;
			ocupation_ne400 : in std_logic;
			correspondence_S123 : in signalStates;
			D07_state : in singleSwitchStates;
			D16_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne992 : in std_logic;
			ocupation_ne994 : in std_logic;
			ocupation_ne993 : in std_logic;
			correspondence_T25 : in signalStates;
			correspondence_J40 : in signalStates;
			Sw05_state : in singleSwitchStates;
			Sw01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_54;
	component railwaySignal_55 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R52_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne123 : in std_logic;
			correspondence_B77 : out signalStates;
			lock_B77 : out objectLock;
			--Ocupation level 1
			ocupation_ne407 : in std_logic;
			ocupation_ne400 : in std_logic;
			correspondence_S123 : in signalStates;
			D07_state : in singleSwitchStates;
			D16_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne992 : in std_logic;
			ocupation_ne994 : in std_logic;
			ocupation_ne993 : in std_logic;
			correspondence_T25 : in signalStates;
			correspondence_J40 : in signalStates;
			Sw05_state : in singleSwitchStates;
			Sw01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_55;
	component railwaySignal_56 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne126 : in std_logic;
			correspondence_T19 : out signalStates;
			lock_T19 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_56;
	component railwaySignal_57 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R14_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne126 : in std_logic;
			correspondence_T20 : out signalStates;
			lock_T20 : out objectLock;
			--Ocupation level 1
			ocupation_ne421 : in std_logic;
			correspondence_T05 : in signalStates;
			D19_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_57;
	component railwaySignal_58 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne127 : in std_logic;
			correspondence_S104 : out signalStates;
			lock_S104 : out objectLock;
			--Ocupation level 1
			ocupation_ne129 : in std_logic;
			ocupation_ne114 : in std_logic;
			ocupation_ne450 : in std_logic;
			correspondence_L29 : in signalStates;
			correspondence_T07 : in signalStates;
			D23_state : in singleSwitchStates;
			D12_state : in doubleSwitchStates;
			correspondence_J48 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_58;
	component railwaySignal_59 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne127 : in std_logic;
			correspondence_S117 : out signalStates;
			lock_S117 : out objectLock;
			--Ocupation level 1
			ocupation_ne135 : in std_logic;
			ocupation_ne910 : in std_logic;
			ocupation_ne101 : in std_logic;
			ocupation_ne134 : in std_logic;
			correspondence_J43 : in signalStates;
			correspondence_T23 : in signalStates;
			D09_state : in singleSwitchStates;
			D10_state : in singleSwitchStates;
			D24_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne100 : in std_logic;
			correspondence_X53 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_59;
	component railwaySignal_60 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R55_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne130 : in std_logic;
			correspondence_C79 : out signalStates;
			lock_C79 : out objectLock;
			--Ocupation level 1
			ocupation_ne910 : in std_logic;
			ocupation_ne101 : in std_logic;
			correspondence_J43 : in signalStates;
			D09_state : in singleSwitchStates;
			D10_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne100 : in std_logic;
			correspondence_X53 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_60;
	component railwaySignal_61 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne130 : in std_logic;
			correspondence_S107 : out signalStates;
			lock_S107 : out objectLock;
			--Ocupation level 1
			ocupation_ne129 : in std_logic;
			ocupation_ne114 : in std_logic;
			ocupation_ne450 : in std_logic;
			correspondence_L29 : in signalStates;
			correspondence_T07 : in signalStates;
			D23_state : in singleSwitchStates;
			D12_state : in doubleSwitchStates;
			correspondence_J48 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_61;
	component railwaySignal_62 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R27_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne132 : in std_logic;
			correspondence_J46 : out signalStates;
			lock_J46 : out objectLock;
			--Ocupation level 1
			ocupation_ne114 : in std_logic;
			correspondence_L29 : in signalStates;
			D23_state : in singleSwitchStates;
			correspondence_J48 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_62;
	component railwaySignal_63 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R28_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne132 : in std_logic;
			correspondence_J47 : out signalStates;
			lock_J47 : out objectLock;
			--Ocupation level 1
			ocupation_ne912 : in std_logic;
			correspondence_J45 : in signalStates;
			D20_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne101 : in std_logic;
			correspondence_J43 : in signalStates;
			D09_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_63;
	component railwaySignal_64 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne133 : in std_logic;
			correspondence_T21 : out signalStates;
			lock_T21 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_64;
	component railwaySignal_65 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R15_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne133 : in std_logic;
			correspondence_T22 : out signalStates;
			lock_T22 : out objectLock;
			--Ocupation level 1
			ocupation_ne465 : in std_logic;
			correspondence_T09 : in signalStates;
			D21_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_65;
	component railwaySignal_66 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne134 : in std_logic;
			correspondence_T23 : out signalStates;
			lock_T23 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_66;
	component railwaySignal_67 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R16_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne134 : in std_logic;
			correspondence_T24 : out signalStates;
			lock_T24 : out objectLock;
			--Ocupation level 1
			ocupation_ne127 : in std_logic;
			correspondence_S104 : in signalStates;
			D24_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne114 : in std_logic;
			ocupation_ne450 : in std_logic;
			ocupation_ne129 : in std_logic;
			correspondence_L29 : in signalStates;
			correspondence_T07 : in signalStates;
			D23_state : in singleSwitchStates;
			D12_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_67;
	component railwaySignal_68 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R56_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne135 : in std_logic;
			correspondence_B80 : out signalStates;
			lock_B80 : out objectLock;
			--Ocupation level 1
			ocupation_ne127 : in std_logic;
			correspondence_S104 : in signalStates;
			D24_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne114 : in std_logic;
			ocupation_ne450 : in std_logic;
			ocupation_ne129 : in std_logic;
			correspondence_L29 : in signalStates;
			correspondence_T07 : in signalStates;
			D23_state : in singleSwitchStates;
			D12_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_68;
	component railwaySignal_69 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R24_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne992 : in std_logic;
			correspondence_J40 : out signalStates;
			lock_J40 : out objectLock;
			--Ocupation level 1
			ocupation_ne100 : in std_logic;
			correspondence_L31 : in signalStates;
			correspondence_X52 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_69;
	component railwaySignal_70 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R80_command : in routeCommands;
			R81_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne992 : in std_logic;
			correspondence_S120 : out signalStates;
			lock_S120 : out objectLock;
			--Ocupation level 1
			ocupation_ne65 : in std_logic;
			ocupation_ne994 : in std_logic;
			ocupation_ne400 : in std_logic;
			correspondence_C94 : in signalStates;
			correspondence_S74 : in signalStates;
			Sw01_state : in singleSwitchStates;
			Sw05_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne63 : in std_logic;
			ocupation_ne407 : in std_logic;
			ocupation_ne404 : in std_logic;
			correspondence_C54 : in signalStates;
			correspondence_C76 : in signalStates;
			correspondence_S93 : in signalStates;
			D18_state : in singleSwitchStates;
			D07_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_70;
	component railwaySignal_71 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne993 : in std_logic;
			correspondence_T25 : out signalStates;
			lock_T25 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_71;
	component railwaySignal_72 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R82_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne993 : in std_logic;
			correspondence_C122 : out signalStates;
			lock_C122 : out objectLock;
			--Ocupation level 1
			ocupation_ne400 : in std_logic;
			correspondence_S74 : in signalStates;
			Sw05_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne407 : in std_logic;
			ocupation_ne404 : in std_logic;
			correspondence_C76 : in signalStates;
			correspondence_S93 : in signalStates;
			D07_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_72;
	component railwaySignal_73 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne995 : in std_logic;
			correspondence_T27 : out signalStates;
			lock_T27 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_73;
	component railwaySignal_74 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R85_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne995 : in std_logic;
			correspondence_C125 : out signalStates;
			lock_C125 : out objectLock;
			--Ocupation level 1
			ocupation_ne297 : in std_logic;
			correspondence_S71 : in signalStates;
			Sw03_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne384 : in std_logic;
			ocupation_ne295 : in std_logic;
			correspondence_C67 : in signalStates;
			correspondence_S84 : in signalStates;
			D04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_74;
	component railwaySignal_75 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R23_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne996 : in std_logic;
			correspondence_J38 : out signalStates;
			lock_J38 : out objectLock;
			--Ocupation level 1
			ocupation_ne98 : in std_logic;
			correspondence_L30 : in signalStates;
			correspondence_X50 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_75;
	component railwaySignal_76 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R88_command : in routeCommands;
			R89_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne996 : in std_logic;
			correspondence_S129 : out signalStates;
			lock_S129 : out objectLock;
			--Ocupation level 1
			ocupation_ne292 : in std_logic;
			ocupation_ne997 : in std_logic;
			ocupation_ne297 : in std_logic;
			correspondence_J37 : in signalStates;
			correspondence_S71 : in signalStates;
			Sw04_state : in singleSwitchStates;
			Sw03_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne290 : in std_logic;
			ocupation_ne384 : in std_logic;
			ocupation_ne295 : in std_logic;
			correspondence_J35 : in signalStates;
			correspondence_C67 : in signalStates;
			correspondence_S84 : in signalStates;
			D14_state : in singleSwitchStates;
			D04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_76;
	component node_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R1_command : in routeCommands;
			R20_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			R41_command : in routeCommands;
			R60_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_0;
	component node_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R35_command : in routeCommands;
			R51_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R64_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_1;
	component node_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			R34_command : in routeCommands;
			R36_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R67_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_2;
	component node_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_3;
	component node_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R38_command : in routeCommands;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			R58_command : in routeCommands;
			R77_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_4;
	component node_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R26_command : in routeCommands;
			R28_command : in routeCommands;
			R37_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_5;
	component node_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R10_command : in routeCommands;
			R17_command : in routeCommands;
			R27_command : in routeCommands;
			R29_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R73_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_6;
	component node_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R39_command : in routeCommands;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			R60_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_7;
	component node_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R2_command : in routeCommands;
			R20_command : in routeCommands;
			R22_command : in routeCommands;
			R40_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_8;
	component node_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R21_command : in routeCommands;
			R22_command : in routeCommands;
			R61_command : in routeCommands;
			R88_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_9;
	component node_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R45_command : in routeCommands;
			R46_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_10;
	component node_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R42_command : in routeCommands;
			R45_command : in routeCommands;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			R87_command : in routeCommands;
			R89_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_11;
	component node_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R2_command : in routeCommands;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			R62_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_12;
	component node_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R42_command : in routeCommands;
			R47_command : in routeCommands;
			R59_command : in routeCommands;
			R60_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_13;
	component node_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R13_command : in routeCommands;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			R52_command : in routeCommands;
			R81_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			R84_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_14;
	component node_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R51_command : in routeCommands;
			R53_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_15;
	component node_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R13_command : in routeCommands;
			R50_command : in routeCommands;
			R52_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_16;
	component node_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			R67_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_17;
	component node_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R7_command : in routeCommands;
			R72_command : in routeCommands;
			R74_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_18;
	component node_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			R75_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_19;
	component node_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R18_command : in routeCommands;
			R23_command : in routeCommands;
			R30_command : in routeCommands;
			R31_command : in routeCommands;
			R34_command : in routeCommands;
			R51_command : in routeCommands;
			R64_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_20;
	component node_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R30_command : in routeCommands;
			R34_command : in routeCommands;
			R35_command : in routeCommands;
			R36_command : in routeCommands;
			R51_command : in routeCommands;
			R64_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_21;
	component node_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R19_command : in routeCommands;
			R24_command : in routeCommands;
			R25_command : in routeCommands;
			R32_command : in routeCommands;
			R33_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_22;
	component node_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			R32_command : in routeCommands;
			R37_command : in routeCommands;
			R38_command : in routeCommands;
			R55_command : in routeCommands;
			R77_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_23;
	component node_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R10_command : in routeCommands;
			R29_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_24;
	component node_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R59_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_25;
	component node_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			R60_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_26;
	component node_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R2_command : in routeCommands;
			R62_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_27;
	component node_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R3_command : in routeCommands;
			R12_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_28;
	component node_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R13_command : in routeCommands;
			R63_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_29;
	component node_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R52_command : in routeCommands;
			R54_command : in routeCommands;
			R64_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_30;
	component node_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			R67_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_31;
	component node_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R5_command : in routeCommands;
			R14_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_32;
	component node_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R16_command : in routeCommands;
			R56_command : in routeCommands;
			R69_command : in routeCommands;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_33;
	component node_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R71_command : in routeCommands;
			R73_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_34;
	component node_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R7_command : in routeCommands;
			R55_command : in routeCommands;
			R57_command : in routeCommands;
			R70_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_35;
	component node_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R75_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_36;
	component node_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R27_command : in routeCommands;
			R28_command : in routeCommands;
			R68_command : in routeCommands;
			R76_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_37;
	component node_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R9_command : in routeCommands;
			R15_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_38;
	component node_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R16_command : in routeCommands;
			R78_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_39;
	component node_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R77_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_40;
	component node_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R24_command : in routeCommands;
			R33_command : in routeCommands;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			R81_command : in routeCommands;
			R84_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_41;
	component node_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_42;
	component node_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R81_command : in routeCommands;
			R84_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_43;
	component node_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_44;
	component node_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R21_command : in routeCommands;
			R23_command : in routeCommands;
			R31_command : in routeCommands;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			R89_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_45;
	component node_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R87_command : in routeCommands;
			R89_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_46;
	component route_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne991_state : in nodeStates;
			ne991_lock : in objectLock;
			ne991_command : out routeCommands;
			T02_state : in signalStates;
			T02_lock : in objectLock;
			T02_command : out routeCommands;
			S64_state : in signalStates;
			routeState : out std_logic
		);
	end component route_0;
	component route_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne377_state : in nodeStates;
			ne377_lock : in objectLock;
			ne377_command : out routeCommands;
			ne111_state : in nodeStates;
			ne111_lock : in objectLock;
			ne111_command : out routeCommands;
			ne290_state : in nodeStates;
			ne290_lock : in objectLock;
			ne290_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_lock : in objectLock;
			D14_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_lock : in objectLock;
			D15_command : out routeCommands;
			T04_state : in signalStates;
			T04_lock : in objectLock;
			T04_command : out routeCommands;
			J35_state : in signalStates;
			routeState : out std_logic
		);
	end component route_1;
	component route_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne377_state : in nodeStates;
			ne377_lock : in objectLock;
			ne377_command : out routeCommands;
			ne113_state : in nodeStates;
			ne113_lock : in objectLock;
			ne113_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_lock : in objectLock;
			D15_command : out routeCommands;
			T04_state : in signalStates;
			T04_lock : in objectLock;
			T04_command : out routeCommands;
			T15_state : in signalStates;
			routeState : out std_logic
		);
	end component route_2;
	component route_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne421_state : in nodeStates;
			ne421_lock : in objectLock;
			ne421_command : out routeCommands;
			ne124_state : in nodeStates;
			ne124_lock : in objectLock;
			ne124_command : out routeCommands;
			ne63_state : in nodeStates;
			ne63_lock : in objectLock;
			ne63_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_lock : in objectLock;
			D18_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_lock : in objectLock;
			D19_command : out routeCommands;
			T06_state : in signalStates;
			T06_lock : in objectLock;
			T06_command : out routeCommands;
			C54_state : in signalStates;
			routeState : out std_logic
		);
	end component route_3;
	component route_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne421_state : in nodeStates;
			ne421_lock : in objectLock;
			ne421_command : out routeCommands;
			ne126_state : in nodeStates;
			ne126_lock : in objectLock;
			ne126_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_lock : in objectLock;
			D19_command : out routeCommands;
			T06_state : in signalStates;
			T06_lock : in objectLock;
			T06_command : out routeCommands;
			T19_state : in signalStates;
			routeState : out std_logic
		);
	end component route_4;
	component route_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne450_state : in nodeStates;
			ne450_lock : in objectLock;
			ne450_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			T08_state : in signalStates;
			T08_lock : in objectLock;
			T08_command : out routeCommands;
			S117_state : in signalStates;
			routeState : out std_logic
		);
	end component route_5;
	component route_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne450_state : in nodeStates;
			ne450_lock : in objectLock;
			ne450_command : out routeCommands;
			ne130_state : in nodeStates;
			ne130_lock : in objectLock;
			ne130_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			T08_state : in signalStates;
			T08_lock : in objectLock;
			T08_command : out routeCommands;
			C79_state : in signalStates;
			routeState : out std_logic
		);
	end component route_6;
	component route_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne465_state : in nodeStates;
			ne465_lock : in objectLock;
			ne465_command : out routeCommands;
			ne131_state : in nodeStates;
			ne131_lock : in objectLock;
			ne131_command : out routeCommands;
			ne912_state : in nodeStates;
			ne912_lock : in objectLock;
			ne912_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_lock : in objectLock;
			D20_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_lock : in objectLock;
			D21_command : out routeCommands;
			T10_state : in signalStates;
			T10_lock : in objectLock;
			T10_command : out routeCommands;
			J45_state : in signalStates;
			routeState : out std_logic
		);
	end component route_7;
	component route_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne465_state : in nodeStates;
			ne465_lock : in objectLock;
			ne465_command : out routeCommands;
			ne133_state : in nodeStates;
			ne133_lock : in objectLock;
			ne133_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_lock : in objectLock;
			D21_command : out routeCommands;
			T10_state : in signalStates;
			T10_lock : in objectLock;
			T10_command : out routeCommands;
			T21_state : in signalStates;
			routeState : out std_logic
		);
	end component route_8;
	component route_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne102_state : in nodeStates;
			ne102_lock : in objectLock;
			ne102_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			T12_state : in signalStates;
			T12_lock : in objectLock;
			T12_command : out routeCommands;
			S101_state : in signalStates;
			routeState : out std_logic
		);
	end component route_9;
	component route_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne104_state : in nodeStates;
			ne104_lock : in objectLock;
			ne104_command : out routeCommands;
			ne384_state : in nodeStates;
			ne384_lock : in objectLock;
			ne384_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_lock : in objectLock;
			D04_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_lock : in objectLock;
			Sw02_command : out routeCommands;
			T14_state : in signalStates;
			T14_lock : in objectLock;
			T14_command : out routeCommands;
			S126_state : in signalStates;
			routeState : out std_logic
		);
	end component route_10;
	component route_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne113_state : in nodeStates;
			ne113_lock : in objectLock;
			ne113_command : out routeCommands;
			ne377_state : in nodeStates;
			ne377_lock : in objectLock;
			ne377_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_lock : in objectLock;
			D15_command : out routeCommands;
			T16_state : in signalStates;
			T16_lock : in objectLock;
			T16_command : out routeCommands;
			T03_state : in signalStates;
			routeState : out std_logic
		);
	end component route_11;
	component route_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne122_state : in nodeStates;
			ne122_lock : in objectLock;
			ne122_command : out routeCommands;
			ne407_state : in nodeStates;
			ne407_lock : in objectLock;
			ne407_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_lock : in objectLock;
			D07_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_lock : in objectLock;
			D16_command : out routeCommands;
			T18_state : in signalStates;
			T18_lock : in objectLock;
			T18_command : out routeCommands;
			S123_state : in signalStates;
			routeState : out std_logic
		);
	end component route_12;
	component route_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne126_state : in nodeStates;
			ne126_lock : in objectLock;
			ne126_command : out routeCommands;
			ne421_state : in nodeStates;
			ne421_lock : in objectLock;
			ne421_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_lock : in objectLock;
			D19_command : out routeCommands;
			T20_state : in signalStates;
			T20_lock : in objectLock;
			T20_command : out routeCommands;
			T05_state : in signalStates;
			routeState : out std_logic
		);
	end component route_13;
	component route_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne133_state : in nodeStates;
			ne133_lock : in objectLock;
			ne133_command : out routeCommands;
			ne465_state : in nodeStates;
			ne465_lock : in objectLock;
			ne465_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_lock : in objectLock;
			D21_command : out routeCommands;
			T22_state : in signalStates;
			T22_lock : in objectLock;
			T22_command : out routeCommands;
			T09_state : in signalStates;
			routeState : out std_logic
		);
	end component route_14;
	component route_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne134_state : in nodeStates;
			ne134_lock : in objectLock;
			ne134_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_lock : in objectLock;
			D24_command : out routeCommands;
			T24_state : in signalStates;
			T24_lock : in objectLock;
			T24_command : out routeCommands;
			S104_state : in signalStates;
			routeState : out std_logic
		);
	end component route_15;
	component route_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			L29_state : in signalStates;
			L29_lock : in objectLock;
			L29_command : out routeCommands;
			J48_state : in signalStates;
			routeState : out std_logic
		);
	end component route_16;
	component route_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			L30_state : in signalStates;
			L30_lock : in objectLock;
			L30_command : out routeCommands;
			X50_state : in signalStates;
			routeState : out std_logic
		);
	end component route_17;
	component route_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			L31_state : in signalStates;
			L31_lock : in objectLock;
			L31_command : out routeCommands;
			X52_state : in signalStates;
			routeState : out std_logic
		);
	end component route_18;
	component route_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne290_state : in nodeStates;
			ne290_lock : in objectLock;
			ne290_command : out routeCommands;
			ne991_state : in nodeStates;
			ne991_lock : in objectLock;
			ne991_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_lock : in objectLock;
			D01_command : out routeCommands;
			J35_state : in signalStates;
			J35_lock : in objectLock;
			J35_command : out routeCommands;
			T01_state : in signalStates;
			routeState : out std_logic
		);
	end component route_19;
	component route_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne292_state : in nodeStates;
			ne292_lock : in objectLock;
			ne292_command : out routeCommands;
			ne996_state : in nodeStates;
			ne996_lock : in objectLock;
			ne996_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			J36_state : in signalStates;
			J36_lock : in objectLock;
			J36_command : out routeCommands;
			J38_state : in signalStates;
			routeState : out std_logic
		);
	end component route_20;
	component route_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne292_state : in nodeStates;
			ne292_lock : in objectLock;
			ne292_command : out routeCommands;
			ne290_state : in nodeStates;
			ne290_lock : in objectLock;
			ne290_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_lock : in objectLock;
			D14_command : out routeCommands;
			J37_state : in signalStates;
			J37_lock : in objectLock;
			J37_command : out routeCommands;
			J35_state : in signalStates;
			routeState : out std_logic
		);
	end component route_21;
	component route_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne996_state : in nodeStates;
			ne996_lock : in objectLock;
			ne996_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			J38_state : in signalStates;
			J38_lock : in objectLock;
			J38_command : out routeCommands;
			L30_state : in signalStates;
			routeState : out std_logic
		);
	end component route_22;
	component route_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne992_state : in nodeStates;
			ne992_lock : in objectLock;
			ne992_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			J40_state : in signalStates;
			J40_lock : in objectLock;
			J40_command : out routeCommands;
			L31_state : in signalStates;
			routeState : out std_logic
		);
	end component route_23;
	component route_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			J43_state : in signalStates;
			J43_lock : in objectLock;
			J43_command : out routeCommands;
			X53_state : in signalStates;
			routeState : out std_logic
		);
	end component route_24;
	component route_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne912_state : in nodeStates;
			ne912_lock : in objectLock;
			ne912_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_lock : in objectLock;
			D09_command : out routeCommands;
			J45_state : in signalStates;
			J45_lock : in objectLock;
			J45_command : out routeCommands;
			J43_state : in signalStates;
			routeState : out std_logic
		);
	end component route_25;
	component route_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne132_state : in nodeStates;
			ne132_lock : in objectLock;
			ne132_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_lock : in objectLock;
			D23_command : out routeCommands;
			J46_state : in signalStates;
			J46_lock : in objectLock;
			J46_command : out routeCommands;
			L29_state : in signalStates;
			routeState : out std_logic
		);
	end component route_26;
	component route_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne132_state : in nodeStates;
			ne132_lock : in objectLock;
			ne132_command : out routeCommands;
			ne912_state : in nodeStates;
			ne912_lock : in objectLock;
			ne912_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_lock : in objectLock;
			D20_command : out routeCommands;
			J47_state : in signalStates;
			J47_lock : in objectLock;
			J47_command : out routeCommands;
			J45_state : in signalStates;
			routeState : out std_logic
		);
	end component route_27;
	component route_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			ne102_state : in nodeStates;
			ne102_lock : in objectLock;
			ne102_command : out routeCommands;
			J48_state : in signalStates;
			J48_lock : in objectLock;
			J48_command : out routeCommands;
			T11_state : in signalStates;
			routeState : out std_logic
		);
	end component route_28;
	component route_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			Lc01_state : in levelCrossingStates;
			Lc01_lock : in objectLock;
			Lc01_command : out routeCommands;
			X50_state : in signalStates;
			X50_lock : in objectLock;
			X50_command : out routeCommands;
			S55_state : in signalStates;
			routeState : out std_logic
		);
	end component route_29;
	component route_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			ne996_state : in nodeStates;
			ne996_lock : in objectLock;
			ne996_command : out routeCommands;
			Lc01_state : in levelCrossingStates;
			Lc01_lock : in objectLock;
			Lc01_command : out routeCommands;
			X51_state : in signalStates;
			X51_lock : in objectLock;
			X51_command : out routeCommands;
			S129_state : in signalStates;
			routeState : out std_logic
		);
	end component route_30;
	component route_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			Lc04_state : in levelCrossingStates;
			Lc04_lock : in objectLock;
			Lc04_command : out routeCommands;
			X52_state : in signalStates;
			X52_lock : in objectLock;
			X52_command : out routeCommands;
			S59_state : in signalStates;
			routeState : out std_logic
		);
	end component route_31;
	component route_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			ne992_state : in nodeStates;
			ne992_lock : in objectLock;
			ne992_command : out routeCommands;
			Lc04_state : in levelCrossingStates;
			Lc04_lock : in objectLock;
			Lc04_command : out routeCommands;
			X53_state : in signalStates;
			X53_lock : in objectLock;
			X53_command : out routeCommands;
			S120_state : in signalStates;
			routeState : out std_logic
		);
	end component route_32;
	component route_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne63_state : in nodeStates;
			ne63_lock : in objectLock;
			ne63_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_lock : in objectLock;
			D05_command : out routeCommands;
			C54_state : in signalStates;
			C54_lock : in objectLock;
			C54_command : out routeCommands;
			X51_state : in signalStates;
			routeState : out std_logic
		);
	end component route_33;
	component route_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			ne61_state : in nodeStates;
			ne61_lock : in objectLock;
			ne61_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_lock : in objectLock;
			D05_command : out routeCommands;
			S55_state : in signalStates;
			S55_lock : in objectLock;
			S55_command : out routeCommands;
			S78_state : in signalStates;
			routeState : out std_logic
		);
	end component route_34;
	component route_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			ne63_state : in nodeStates;
			ne63_lock : in objectLock;
			ne63_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_lock : in objectLock;
			D05_command : out routeCommands;
			S55_state : in signalStates;
			S55_lock : in objectLock;
			S55_command : out routeCommands;
			S95_state : in signalStates;
			routeState : out std_logic
		);
	end component route_35;
	component route_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			ne912_state : in nodeStates;
			ne912_lock : in objectLock;
			ne912_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_lock : in objectLock;
			D09_command : out routeCommands;
			S59_state : in signalStates;
			S59_lock : in objectLock;
			S59_command : out routeCommands;
			S110_state : in signalStates;
			routeState : out std_logic
		);
	end component route_36;
	component route_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			ne910_state : in nodeStates;
			ne910_lock : in objectLock;
			ne910_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_lock : in objectLock;
			D09_command : out routeCommands;
			S59_state : in signalStates;
			S59_lock : in objectLock;
			S59_command : out routeCommands;
			S81_state : in signalStates;
			routeState : out std_logic
		);
	end component route_37;
	component route_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne991_state : in nodeStates;
			ne991_lock : in objectLock;
			ne991_command : out routeCommands;
			ne288_state : in nodeStates;
			ne288_lock : in objectLock;
			ne288_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_lock : in objectLock;
			D01_command : out routeCommands;
			S64_state : in signalStates;
			S64_lock : in objectLock;
			S64_command : out routeCommands;
			S69_state : in signalStates;
			routeState : out std_logic
		);
	end component route_38;
	component route_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne991_state : in nodeStates;
			ne991_lock : in objectLock;
			ne991_command : out routeCommands;
			ne290_state : in nodeStates;
			ne290_lock : in objectLock;
			ne290_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_lock : in objectLock;
			D01_command : out routeCommands;
			S64_state : in signalStates;
			S64_lock : in objectLock;
			S64_command : out routeCommands;
			S86_state : in signalStates;
			routeState : out std_logic
		);
	end component route_39;
	component route_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne295_state : in nodeStates;
			ne295_lock : in objectLock;
			ne295_command : out routeCommands;
			ne288_state : in nodeStates;
			ne288_lock : in objectLock;
			ne288_command : out routeCommands;
			ne991_state : in nodeStates;
			ne991_lock : in objectLock;
			ne991_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_lock : in objectLock;
			D01_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_lock : in objectLock;
			D03_command : out routeCommands;
			C67_state : in signalStates;
			C67_lock : in objectLock;
			C67_command : out routeCommands;
			T01_state : in signalStates;
			routeState : out std_logic
		);
	end component route_40;
	component route_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			ne384_state : in nodeStates;
			ne384_lock : in objectLock;
			ne384_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_lock : in objectLock;
			D04_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_lock : in objectLock;
			Sw02_command : out routeCommands;
			B68_state : in signalStates;
			B68_lock : in objectLock;
			B68_command : out routeCommands;
			S126_state : in signalStates;
			routeState : out std_logic
		);
	end component route_41;
	component route_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne288_state : in nodeStates;
			ne288_lock : in objectLock;
			ne288_command : out routeCommands;
			ne295_state : in nodeStates;
			ne295_lock : in objectLock;
			ne295_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_lock : in objectLock;
			D03_command : out routeCommands;
			S69_state : in signalStates;
			S69_lock : in objectLock;
			S69_command : out routeCommands;
			C70_state : in signalStates;
			routeState : out std_logic
		);
	end component route_42;
	component route_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne288_state : in nodeStates;
			ne288_lock : in objectLock;
			ne288_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_lock : in objectLock;
			D03_command : out routeCommands;
			S69_state : in signalStates;
			S69_lock : in objectLock;
			S69_command : out routeCommands;
			B68_state : in signalStates;
			routeState : out std_logic
		);
	end component route_43;
	component route_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne295_state : in nodeStates;
			ne295_lock : in objectLock;
			ne295_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_lock : in objectLock;
			D04_command : out routeCommands;
			C70_state : in signalStates;
			C70_lock : in objectLock;
			C70_command : out routeCommands;
			S126_state : in signalStates;
			routeState : out std_logic
		);
	end component route_44;
	component route_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			ne295_state : in nodeStates;
			ne295_lock : in objectLock;
			ne295_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_lock : in objectLock;
			D04_command : out routeCommands;
			S71_state : in signalStates;
			S71_lock : in objectLock;
			S71_command : out routeCommands;
			C67_state : in signalStates;
			routeState : out std_logic
		);
	end component route_45;
	component route_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			ne384_state : in nodeStates;
			ne384_lock : in objectLock;
			ne384_command : out routeCommands;
			D04_state : in singleSwitchStates;
			D04_lock : in objectLock;
			D04_command : out routeCommands;
			S71_state : in signalStates;
			S71_lock : in objectLock;
			S71_command : out routeCommands;
			S84_state : in signalStates;
			routeState : out std_logic
		);
	end component route_46;
	component route_47 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne404_state : in nodeStates;
			ne404_lock : in objectLock;
			ne404_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_lock : in objectLock;
			D07_command : out routeCommands;
			C73_state : in signalStates;
			C73_lock : in objectLock;
			C73_command : out routeCommands;
			S123_state : in signalStates;
			routeState : out std_logic
		);
	end component route_47;
	component route_48 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			ne404_state : in nodeStates;
			ne404_lock : in objectLock;
			ne404_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_lock : in objectLock;
			D07_command : out routeCommands;
			S74_state : in signalStates;
			S74_lock : in objectLock;
			S74_command : out routeCommands;
			C76_state : in signalStates;
			routeState : out std_logic
		);
	end component route_48;
	component route_49 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			ne407_state : in nodeStates;
			ne407_lock : in objectLock;
			ne407_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_lock : in objectLock;
			D07_command : out routeCommands;
			S74_state : in signalStates;
			S74_lock : in objectLock;
			S74_command : out routeCommands;
			S93_state : in signalStates;
			routeState : out std_logic
		);
	end component route_49;
	component route_50 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne404_state : in nodeStates;
			ne404_lock : in objectLock;
			ne404_command : out routeCommands;
			ne61_state : in nodeStates;
			ne61_lock : in objectLock;
			ne61_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_lock : in objectLock;
			D05_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_lock : in objectLock;
			D08_command : out routeCommands;
			C76_state : in signalStates;
			C76_lock : in objectLock;
			C76_command : out routeCommands;
			X51_state : in signalStates;
			routeState : out std_logic
		);
	end component route_50;
	component route_51 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne123_state : in nodeStates;
			ne123_lock : in objectLock;
			ne123_command : out routeCommands;
			ne407_state : in nodeStates;
			ne407_lock : in objectLock;
			ne407_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			D07_state : in singleSwitchStates;
			D07_lock : in objectLock;
			D07_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_lock : in objectLock;
			D16_command : out routeCommands;
			B77_state : in signalStates;
			B77_lock : in objectLock;
			B77_command : out routeCommands;
			S123_state : in signalStates;
			routeState : out std_logic
		);
	end component route_51;
	component route_52 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne61_state : in nodeStates;
			ne61_lock : in objectLock;
			ne61_command : out routeCommands;
			ne404_state : in nodeStates;
			ne404_lock : in objectLock;
			ne404_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_lock : in objectLock;
			D08_command : out routeCommands;
			S78_state : in signalStates;
			S78_lock : in objectLock;
			S78_command : out routeCommands;
			C73_state : in signalStates;
			routeState : out std_logic
		);
	end component route_52;
	component route_53 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne61_state : in nodeStates;
			ne61_lock : in objectLock;
			ne61_command : out routeCommands;
			ne123_state : in nodeStates;
			ne123_lock : in objectLock;
			ne123_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_lock : in objectLock;
			D08_command : out routeCommands;
			S78_state : in signalStates;
			S78_lock : in objectLock;
			S78_command : out routeCommands;
			B77_state : in signalStates;
			routeState : out std_logic
		);
	end component route_53;
	component route_54 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne130_state : in nodeStates;
			ne130_lock : in objectLock;
			ne130_command : out routeCommands;
			ne910_state : in nodeStates;
			ne910_lock : in objectLock;
			ne910_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_lock : in objectLock;
			D09_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_lock : in objectLock;
			D10_command : out routeCommands;
			C79_state : in signalStates;
			C79_lock : in objectLock;
			C79_command : out routeCommands;
			J43_state : in signalStates;
			routeState : out std_logic
		);
	end component route_54;
	component route_55 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne135_state : in nodeStates;
			ne135_lock : in objectLock;
			ne135_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_lock : in objectLock;
			D24_command : out routeCommands;
			B80_state : in signalStates;
			B80_lock : in objectLock;
			B80_command : out routeCommands;
			S104_state : in signalStates;
			routeState : out std_logic
		);
	end component route_55;
	component route_56 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne910_state : in nodeStates;
			ne910_lock : in objectLock;
			ne910_command : out routeCommands;
			ne130_state : in nodeStates;
			ne130_lock : in objectLock;
			ne130_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_lock : in objectLock;
			D10_command : out routeCommands;
			S81_state : in signalStates;
			S81_lock : in objectLock;
			S81_command : out routeCommands;
			S107_state : in signalStates;
			routeState : out std_logic
		);
	end component route_56;
	component route_57 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne910_state : in nodeStates;
			ne910_lock : in objectLock;
			ne910_command : out routeCommands;
			ne135_state : in nodeStates;
			ne135_lock : in objectLock;
			ne135_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_lock : in objectLock;
			D10_command : out routeCommands;
			S81_state : in signalStates;
			S81_lock : in objectLock;
			S81_command : out routeCommands;
			B80_state : in signalStates;
			routeState : out std_logic
		);
	end component route_57;
	component route_58 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne384_state : in nodeStates;
			ne384_lock : in objectLock;
			ne384_command : out routeCommands;
			ne104_state : in nodeStates;
			ne104_lock : in objectLock;
			ne104_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_lock : in objectLock;
			Sw02_command : out routeCommands;
			S84_state : in signalStates;
			S84_lock : in objectLock;
			S84_command : out routeCommands;
			T13_state : in signalStates;
			routeState : out std_logic
		);
	end component route_58;
	component route_59 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne384_state : in nodeStates;
			ne384_lock : in objectLock;
			ne384_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			ne288_state : in nodeStates;
			ne288_lock : in objectLock;
			ne288_command : out routeCommands;
			ne991_state : in nodeStates;
			ne991_lock : in objectLock;
			ne991_command : out routeCommands;
			D01_state : in singleSwitchStates;
			D01_lock : in objectLock;
			D01_command : out routeCommands;
			D03_state : in singleSwitchStates;
			D03_lock : in objectLock;
			D03_command : out routeCommands;
			Sw02_state : in singleSwitchStates;
			Sw02_lock : in objectLock;
			Sw02_command : out routeCommands;
			S84_state : in signalStates;
			S84_lock : in objectLock;
			S84_command : out routeCommands;
			T01_state : in signalStates;
			routeState : out std_logic
		);
	end component route_59;
	component route_60 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne290_state : in nodeStates;
			ne290_lock : in objectLock;
			ne290_command : out routeCommands;
			ne292_state : in nodeStates;
			ne292_lock : in objectLock;
			ne292_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_lock : in objectLock;
			D14_command : out routeCommands;
			S86_state : in signalStates;
			S86_lock : in objectLock;
			S86_command : out routeCommands;
			J36_state : in signalStates;
			routeState : out std_logic
		);
	end component route_60;
	component route_61 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne290_state : in nodeStates;
			ne290_lock : in objectLock;
			ne290_command : out routeCommands;
			ne111_state : in nodeStates;
			ne111_lock : in objectLock;
			ne111_command : out routeCommands;
			ne377_state : in nodeStates;
			ne377_lock : in objectLock;
			ne377_command : out routeCommands;
			D14_state : in singleSwitchStates;
			D14_lock : in objectLock;
			D14_command : out routeCommands;
			D15_state : in singleSwitchStates;
			D15_lock : in objectLock;
			D15_command : out routeCommands;
			S86_state : in signalStates;
			S86_lock : in objectLock;
			S86_command : out routeCommands;
			T03_state : in signalStates;
			routeState : out std_logic
		);
	end component route_61;
	component route_62 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne407_state : in nodeStates;
			ne407_lock : in objectLock;
			ne407_command : out routeCommands;
			ne122_state : in nodeStates;
			ne122_lock : in objectLock;
			ne122_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_lock : in objectLock;
			D16_command : out routeCommands;
			S93_state : in signalStates;
			S93_lock : in objectLock;
			S93_command : out routeCommands;
			T17_state : in signalStates;
			routeState : out std_logic
		);
	end component route_62;
	component route_63 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne407_state : in nodeStates;
			ne407_lock : in objectLock;
			ne407_command : out routeCommands;
			ne123_state : in nodeStates;
			ne123_lock : in objectLock;
			ne123_command : out routeCommands;
			ne61_state : in nodeStates;
			ne61_lock : in objectLock;
			ne61_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			D05_state : in singleSwitchStates;
			D05_lock : in objectLock;
			D05_command : out routeCommands;
			D08_state : in singleSwitchStates;
			D08_lock : in objectLock;
			D08_command : out routeCommands;
			D16_state : in singleSwitchStates;
			D16_lock : in objectLock;
			D16_command : out routeCommands;
			S93_state : in signalStates;
			S93_lock : in objectLock;
			S93_command : out routeCommands;
			X51_state : in signalStates;
			routeState : out std_logic
		);
	end component route_63;
	component route_64 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne65_state : in nodeStates;
			ne65_lock : in objectLock;
			ne65_command : out routeCommands;
			ne63_state : in nodeStates;
			ne63_lock : in objectLock;
			ne63_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_lock : in objectLock;
			D18_command : out routeCommands;
			C94_state : in signalStates;
			C94_lock : in objectLock;
			C94_command : out routeCommands;
			C54_state : in signalStates;
			routeState : out std_logic
		);
	end component route_64;
	component route_65 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne63_state : in nodeStates;
			ne63_lock : in objectLock;
			ne63_command : out routeCommands;
			ne65_state : in nodeStates;
			ne65_lock : in objectLock;
			ne65_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_lock : in objectLock;
			D18_command : out routeCommands;
			S95_state : in signalStates;
			S95_lock : in objectLock;
			S95_command : out routeCommands;
			C119_state : in signalStates;
			routeState : out std_logic
		);
	end component route_65;
	component route_66 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne63_state : in nodeStates;
			ne63_lock : in objectLock;
			ne63_command : out routeCommands;
			ne124_state : in nodeStates;
			ne124_lock : in objectLock;
			ne124_command : out routeCommands;
			ne421_state : in nodeStates;
			ne421_lock : in objectLock;
			ne421_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_lock : in objectLock;
			D18_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_lock : in objectLock;
			D19_command : out routeCommands;
			S95_state : in signalStates;
			S95_lock : in objectLock;
			S95_command : out routeCommands;
			T05_state : in signalStates;
			routeState : out std_logic
		);
	end component route_66;
	component route_67 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			ne132_state : in nodeStates;
			ne132_lock : in objectLock;
			ne132_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_lock : in objectLock;
			D23_command : out routeCommands;
			S101_state : in signalStates;
			S101_lock : in objectLock;
			S101_command : out routeCommands;
			J47_state : in signalStates;
			routeState : out std_logic
		);
	end component route_67;
	component route_68 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_lock : in objectLock;
			ne129_command : out routeCommands;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_lock : in objectLock;
			D23_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			S101_state : in signalStates;
			S101_lock : in objectLock;
			S101_command : out routeCommands;
			S117_state : in signalStates;
			routeState : out std_logic
		);
	end component route_68;
	component route_69 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_lock : in objectLock;
			ne129_command : out routeCommands;
			ne130_state : in nodeStates;
			ne130_lock : in objectLock;
			ne130_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_lock : in objectLock;
			D23_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			S101_state : in signalStates;
			S101_lock : in objectLock;
			S101_command : out routeCommands;
			C79_state : in signalStates;
			routeState : out std_logic
		);
	end component route_69;
	component route_70 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_lock : in objectLock;
			ne129_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_lock : in objectLock;
			D23_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			S104_state : in signalStates;
			S104_lock : in objectLock;
			S104_command : out routeCommands;
			L29_state : in signalStates;
			routeState : out std_logic
		);
	end component route_70;
	component route_71 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			ne450_state : in nodeStates;
			ne450_lock : in objectLock;
			ne450_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			S104_state : in signalStates;
			S104_lock : in objectLock;
			S104_command : out routeCommands;
			T07_state : in signalStates;
			routeState : out std_logic
		);
	end component route_71;
	component route_72 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne130_state : in nodeStates;
			ne130_lock : in objectLock;
			ne130_command : out routeCommands;
			ne129_state : in nodeStates;
			ne129_lock : in objectLock;
			ne129_command : out routeCommands;
			ne114_state : in nodeStates;
			ne114_lock : in objectLock;
			ne114_command : out routeCommands;
			D23_state : in singleSwitchStates;
			D23_lock : in objectLock;
			D23_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			S107_state : in signalStates;
			S107_lock : in objectLock;
			S107_command : out routeCommands;
			L29_state : in signalStates;
			routeState : out std_logic
		);
	end component route_72;
	component route_73 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne130_state : in nodeStates;
			ne130_lock : in objectLock;
			ne130_command : out routeCommands;
			ne450_state : in nodeStates;
			ne450_lock : in objectLock;
			ne450_command : out routeCommands;
			D12_state : in doubleSwitchStates;
			D12_lock : in objectLock;
			D12_command : out routeCommands;
			S107_state : in signalStates;
			S107_lock : in objectLock;
			S107_command : out routeCommands;
			T07_state : in signalStates;
			routeState : out std_logic
		);
	end component route_73;
	component route_74 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne912_state : in nodeStates;
			ne912_lock : in objectLock;
			ne912_command : out routeCommands;
			ne131_state : in nodeStates;
			ne131_lock : in objectLock;
			ne131_command : out routeCommands;
			ne465_state : in nodeStates;
			ne465_lock : in objectLock;
			ne465_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_lock : in objectLock;
			D20_command : out routeCommands;
			D21_state : in singleSwitchStates;
			D21_lock : in objectLock;
			D21_command : out routeCommands;
			S110_state : in signalStates;
			S110_lock : in objectLock;
			S110_command : out routeCommands;
			T09_state : in signalStates;
			routeState : out std_logic
		);
	end component route_74;
	component route_75 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne912_state : in nodeStates;
			ne912_lock : in objectLock;
			ne912_command : out routeCommands;
			ne132_state : in nodeStates;
			ne132_lock : in objectLock;
			ne132_command : out routeCommands;
			D20_state : in singleSwitchStates;
			D20_lock : in objectLock;
			D20_command : out routeCommands;
			S110_state : in signalStates;
			S110_lock : in objectLock;
			S110_command : out routeCommands;
			J46_state : in signalStates;
			routeState : out std_logic
		);
	end component route_75;
	component route_76 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			ne135_state : in nodeStates;
			ne135_lock : in objectLock;
			ne135_command : out routeCommands;
			ne910_state : in nodeStates;
			ne910_lock : in objectLock;
			ne910_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			D09_state : in singleSwitchStates;
			D09_lock : in objectLock;
			D09_command : out routeCommands;
			D10_state : in singleSwitchStates;
			D10_lock : in objectLock;
			D10_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_lock : in objectLock;
			D24_command : out routeCommands;
			S117_state : in signalStates;
			S117_lock : in objectLock;
			S117_command : out routeCommands;
			J43_state : in signalStates;
			routeState : out std_logic
		);
	end component route_76;
	component route_77 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne127_state : in nodeStates;
			ne127_lock : in objectLock;
			ne127_command : out routeCommands;
			ne134_state : in nodeStates;
			ne134_lock : in objectLock;
			ne134_command : out routeCommands;
			D24_state : in singleSwitchStates;
			D24_lock : in objectLock;
			D24_command : out routeCommands;
			S117_state : in signalStates;
			S117_lock : in objectLock;
			S117_command : out routeCommands;
			T23_state : in signalStates;
			routeState : out std_logic
		);
	end component route_77;
	component route_78 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne65_state : in nodeStates;
			ne65_lock : in objectLock;
			ne65_command : out routeCommands;
			ne992_state : in nodeStates;
			ne992_lock : in objectLock;
			ne992_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_lock : in objectLock;
			Sw01_command : out routeCommands;
			C119_state : in signalStates;
			C119_lock : in objectLock;
			C119_command : out routeCommands;
			J40_state : in signalStates;
			routeState : out std_logic
		);
	end component route_78;
	component route_79 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne992_state : in nodeStates;
			ne992_lock : in objectLock;
			ne992_command : out routeCommands;
			ne65_state : in nodeStates;
			ne65_lock : in objectLock;
			ne65_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_lock : in objectLock;
			Sw01_command : out routeCommands;
			S120_state : in signalStates;
			S120_lock : in objectLock;
			S120_command : out routeCommands;
			C94_state : in signalStates;
			routeState : out std_logic
		);
	end component route_79;
	component route_80 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne992_state : in nodeStates;
			ne992_lock : in objectLock;
			ne992_command : out routeCommands;
			ne994_state : in nodeStates;
			ne994_lock : in objectLock;
			ne994_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_lock : in objectLock;
			Sw01_command : out routeCommands;
			Sw05_state : in singleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			S120_state : in signalStates;
			S120_lock : in objectLock;
			S120_command : out routeCommands;
			S74_state : in signalStates;
			routeState : out std_logic
		);
	end component route_80;
	component route_81 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne993_state : in nodeStates;
			ne993_lock : in objectLock;
			ne993_command : out routeCommands;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			Sw05_state : in singleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			C122_state : in signalStates;
			C122_lock : in objectLock;
			C122_command : out routeCommands;
			S74_state : in signalStates;
			routeState : out std_logic
		);
	end component route_81;
	component route_82 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			ne993_state : in nodeStates;
			ne993_lock : in objectLock;
			ne993_command : out routeCommands;
			Sw05_state : in singleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			S123_state : in signalStates;
			S123_lock : in objectLock;
			S123_command : out routeCommands;
			T25_state : in signalStates;
			routeState : out std_logic
		);
	end component route_82;
	component route_83 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne400_state : in nodeStates;
			ne400_lock : in objectLock;
			ne400_command : out routeCommands;
			ne994_state : in nodeStates;
			ne994_lock : in objectLock;
			ne994_command : out routeCommands;
			ne992_state : in nodeStates;
			ne992_lock : in objectLock;
			ne992_command : out routeCommands;
			Sw01_state : in singleSwitchStates;
			Sw01_lock : in objectLock;
			Sw01_command : out routeCommands;
			Sw05_state : in singleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			S123_state : in signalStates;
			S123_lock : in objectLock;
			S123_command : out routeCommands;
			J40_state : in signalStates;
			routeState : out std_logic
		);
	end component route_83;
	component route_84 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne995_state : in nodeStates;
			ne995_lock : in objectLock;
			ne995_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			C125_state : in signalStates;
			C125_lock : in objectLock;
			C125_command : out routeCommands;
			S71_state : in signalStates;
			routeState : out std_logic
		);
	end component route_84;
	component route_85 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			ne995_state : in nodeStates;
			ne995_lock : in objectLock;
			ne995_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			S126_state : in signalStates;
			S126_lock : in objectLock;
			S126_command : out routeCommands;
			T27_state : in signalStates;
			routeState : out std_logic
		);
	end component route_85;
	component route_86 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			ne997_state : in nodeStates;
			ne997_lock : in objectLock;
			ne997_command : out routeCommands;
			ne996_state : in nodeStates;
			ne996_lock : in objectLock;
			ne996_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			S126_state : in signalStates;
			S126_lock : in objectLock;
			S126_command : out routeCommands;
			J38_state : in signalStates;
			routeState : out std_logic
		);
	end component route_86;
	component route_87 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne996_state : in nodeStates;
			ne996_lock : in objectLock;
			ne996_command : out routeCommands;
			ne292_state : in nodeStates;
			ne292_lock : in objectLock;
			ne292_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			S129_state : in signalStates;
			S129_lock : in objectLock;
			S129_command : out routeCommands;
			J37_state : in signalStates;
			routeState : out std_logic
		);
	end component route_87;
	component route_88 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne996_state : in nodeStates;
			ne996_lock : in objectLock;
			ne996_command : out routeCommands;
			ne997_state : in nodeStates;
			ne997_lock : in objectLock;
			ne997_command : out routeCommands;
			ne297_state : in nodeStates;
			ne297_lock : in objectLock;
			ne297_command : out routeCommands;
			Sw03_state : in singleSwitchStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			S129_state : in signalStates;
			S129_lock : in objectLock;
			S129_command : out routeCommands;
			S71_state : in signalStates;
			routeState : out std_logic
		);
	end component route_88;
	signal state_Lc01 , state_Lc04 : levelCrossingStates;
	signal Lc01_locking , Lc04_locking : objectLock;
	signal state_D01 , state_D08 , state_D05 , state_D18 , state_Sw01 , state_D10 , state_D09 , state_D20 , state_D23 , state_D03 , state_D14 , state_Sw04 , state_D04 , state_Sw03 , state_D15 , state_Sw02 , state_D07 , state_Sw05 , state_D16 , state_D19 , state_D21 , state_D24 : singleSwitchStates;
	signal D01_locking , D08_locking , D05_locking , D18_locking , Sw01_locking , D10_locking , D09_locking , D20_locking , D23_locking , D03_locking , D14_locking , Sw04_locking , D04_locking , Sw03_locking , D15_locking , Sw02_locking , D07_locking , Sw05_locking , D16_locking , D19_locking , D21_locking , D24_locking : objectLock;
	signal state_D12 : doubleSwitchStates;
	signal D12_locking : objectLock;
	signal state_T01 , state_T02 , state_S64 , state_S78 , state_C54 , state_S95 , state_C94 , state_C119 , state_S81 , state_J45 , state_S110 , state_L29 , state_J48 , state_S101 , state_S69 , state_J35 , state_S86 , state_J36 , state_J37 , state_C67 , state_C70 , state_S71 , state_S126 , state_T03 , state_T04 , state_S84 , state_S74 , state_S123 , state_C73 , state_C76 , state_S93 , state_T05 , state_T06 , state_T07 , state_T08 , state_T09 , state_T10 , state_L30 , state_X50 , state_X51 , state_S55 , state_L31 , state_X52 , state_X53 , state_J43 , state_S59 , state_T11 , state_T12 , state_T13 , state_T14 , state_B68 , state_T15 , state_T16 , state_T17 , state_T18 , state_B77 , state_T19 , state_T20 , state_S104 , state_S117 , state_C79 , state_S107 , state_J46 , state_J47 , state_T21 , state_T22 , state_T23 , state_T24 , state_B80 , state_J40 , state_S120 , state_T25 , state_C122 , state_T27 , state_C125 , state_J38 , state_S129 : signalStates;
	signal T01_locking , T02_locking , S64_locking , S78_locking , C54_locking , S95_locking , C94_locking , C119_locking , S81_locking , J45_locking , S110_locking , L29_locking , J48_locking , S101_locking , S69_locking , J35_locking , S86_locking , J36_locking , J37_locking , C67_locking , C70_locking , S71_locking , S126_locking , T03_locking , T04_locking , S84_locking , S74_locking , S123_locking , C73_locking , C76_locking , S93_locking , T05_locking , T06_locking , T07_locking , T08_locking , T09_locking , T10_locking , L30_locking , X50_locking , X51_locking , S55_locking , L31_locking , X52_locking , X53_locking , J43_locking , S59_locking , T11_locking , T12_locking , T13_locking , T14_locking , B68_locking , T15_locking , T16_locking , T17_locking , T18_locking , B77_locking , T19_locking , T20_locking , S104_locking , S117_locking , C79_locking , S107_locking , J46_locking , J47_locking , T21_locking , T22_locking , T23_locking , T24_locking , B80_locking , J40_locking , S120_locking , T25_locking , C122_locking , T27_locking , C125_locking , J38_locking , S129_locking : objectLock;
	signal state_ne991 , state_ne61 , state_ne63 , state_ne65 , state_ne910 , state_ne912 , state_ne114 , state_ne288 , state_ne290 , state_ne292 , state_ne295 , state_ne297 , state_ne377 , state_ne384 , state_ne400 , state_ne404 , state_ne407 , state_ne421 , state_ne450 , state_ne465 , state_ne98 , state_ne99 , state_ne100 , state_ne101 , state_ne102 , state_ne104 , state_ne110 , state_ne111 , state_ne113 , state_ne122 , state_ne123 , state_ne124 , state_ne126 , state_ne127 , state_ne129 , state_ne130 , state_ne131 , state_ne132 , state_ne133 , state_ne134 , state_ne135 , state_ne992 , state_ne993 , state_ne994 , state_ne995 , state_ne996 , state_ne997 : nodeStates;
	signal ne991_locking , ne61_locking , ne63_locking , ne65_locking , ne910_locking , ne912_locking , ne114_locking , ne288_locking , ne290_locking , ne292_locking , ne295_locking , ne297_locking , ne377_locking , ne384_locking , ne400_locking , ne404_locking , ne407_locking , ne421_locking , ne450_locking , ne465_locking , ne98_locking , ne99_locking , ne100_locking , ne101_locking , ne102_locking , ne104_locking , ne110_locking , ne111_locking , ne113_locking , ne122_locking , ne123_locking , ne124_locking , ne126_locking , ne127_locking , ne129_locking , ne130_locking , ne131_locking , ne132_locking , ne133_locking , ne134_locking , ne135_locking , ne992_locking , ne993_locking , ne994_locking , ne995_locking , ne996_locking , ne997_locking : objectLock;
	signal cmd_R1_ne991 , cmd_R2_ne377 , cmd_R2_ne111 , cmd_R2_ne290 , cmd_R3_ne377 , cmd_R3_ne113 , cmd_R4_ne421 , cmd_R4_ne124 , cmd_R4_ne63 , cmd_R5_ne421 , cmd_R5_ne126 , cmd_R6_ne450 , cmd_R6_ne127 , cmd_R7_ne450 , cmd_R7_ne130 , cmd_R8_ne465 , cmd_R8_ne131 , cmd_R8_ne912 , cmd_R9_ne465 , cmd_R9_ne133 , cmd_R10_ne102 , cmd_R10_ne114 , cmd_R11_ne104 , cmd_R11_ne384 , cmd_R11_ne297 , cmd_R12_ne113 , cmd_R12_ne377 , cmd_R13_ne122 , cmd_R13_ne407 , cmd_R13_ne400 , cmd_R14_ne126 , cmd_R14_ne421 , cmd_R15_ne133 , cmd_R15_ne465 , cmd_R16_ne134 , cmd_R16_ne127 , cmd_R17_ne114 , cmd_R18_ne98 , cmd_R19_ne100 , cmd_R20_ne290 , cmd_R20_ne991 , cmd_R21_ne292 , cmd_R21_ne996 , cmd_R22_ne292 , cmd_R22_ne290 , cmd_R23_ne996 , cmd_R23_ne98 , cmd_R24_ne992 , cmd_R24_ne100 , cmd_R25_ne101 , cmd_R25_ne100 , cmd_R26_ne912 , cmd_R26_ne101 , cmd_R27_ne132 , cmd_R27_ne114 , cmd_R28_ne132 , cmd_R28_ne912 , cmd_R29_ne114 , cmd_R29_ne102 , cmd_R30_ne98 , cmd_R30_ne99 , cmd_R31_ne98 , cmd_R31_ne996 , cmd_R32_ne100 , cmd_R32_ne101 , cmd_R33_ne100 , cmd_R33_ne992 , cmd_R34_ne63 , cmd_R34_ne99 , cmd_R34_ne98 , cmd_R35_ne99 , cmd_R35_ne61 , cmd_R36_ne99 , cmd_R36_ne63 , cmd_R37_ne101 , cmd_R37_ne912 , cmd_R38_ne101 , cmd_R38_ne910 , cmd_R39_ne991 , cmd_R39_ne288 , cmd_R40_ne991 , cmd_R40_ne290 , cmd_R41_ne295 , cmd_R41_ne288 , cmd_R41_ne991 , cmd_R42_ne110 , cmd_R42_ne384 , cmd_R42_ne297 , cmd_R43_ne288 , cmd_R43_ne295 , cmd_R44_ne288 , cmd_R44_ne110 , cmd_R45_ne295 , cmd_R45_ne297 , cmd_R46_ne297 , cmd_R46_ne295 , cmd_R47_ne297 , cmd_R47_ne384 , cmd_R48_ne404 , cmd_R48_ne400 , cmd_R49_ne400 , cmd_R49_ne404 , cmd_R50_ne400 , cmd_R50_ne407 , cmd_R51_ne404 , cmd_R51_ne61 , cmd_R51_ne99 , cmd_R51_ne98 , cmd_R52_ne123 , cmd_R52_ne407 , cmd_R52_ne400 , cmd_R53_ne61 , cmd_R53_ne404 , cmd_R54_ne61 , cmd_R54_ne123 , cmd_R55_ne130 , cmd_R55_ne910 , cmd_R55_ne101 , cmd_R56_ne135 , cmd_R56_ne127 , cmd_R57_ne910 , cmd_R57_ne130 , cmd_R58_ne910 , cmd_R58_ne135 , cmd_R59_ne384 , cmd_R59_ne104 , cmd_R60_ne384 , cmd_R60_ne110 , cmd_R60_ne288 , cmd_R60_ne991 , cmd_R61_ne290 , cmd_R61_ne292 , cmd_R62_ne290 , cmd_R62_ne111 , cmd_R62_ne377 , cmd_R63_ne407 , cmd_R63_ne122 , cmd_R64_ne407 , cmd_R64_ne123 , cmd_R64_ne61 , cmd_R64_ne99 , cmd_R64_ne98 , cmd_R65_ne65 , cmd_R65_ne63 , cmd_R66_ne63 , cmd_R66_ne65 , cmd_R67_ne63 , cmd_R67_ne124 , cmd_R67_ne421 , cmd_R68_ne114 , cmd_R68_ne132 , cmd_R69_ne114 , cmd_R69_ne129 , cmd_R69_ne127 , cmd_R70_ne114 , cmd_R70_ne129 , cmd_R70_ne130 , cmd_R71_ne127 , cmd_R71_ne129 , cmd_R71_ne114 , cmd_R72_ne127 , cmd_R72_ne450 , cmd_R73_ne130 , cmd_R73_ne129 , cmd_R73_ne114 , cmd_R74_ne130 , cmd_R74_ne450 , cmd_R75_ne912 , cmd_R75_ne131 , cmd_R75_ne465 , cmd_R76_ne912 , cmd_R76_ne132 , cmd_R77_ne127 , cmd_R77_ne135 , cmd_R77_ne910 , cmd_R77_ne101 , cmd_R78_ne127 , cmd_R78_ne134 , cmd_R79_ne65 , cmd_R79_ne992 , cmd_R80_ne992 , cmd_R80_ne65 , cmd_R81_ne992 , cmd_R81_ne994 , cmd_R81_ne400 , cmd_R82_ne993 , cmd_R82_ne400 , cmd_R83_ne400 , cmd_R83_ne993 , cmd_R84_ne400 , cmd_R84_ne994 , cmd_R84_ne992 , cmd_R85_ne995 , cmd_R85_ne297 , cmd_R86_ne297 , cmd_R86_ne995 , cmd_R87_ne297 , cmd_R87_ne997 , cmd_R87_ne996 , cmd_R88_ne996 , cmd_R88_ne292 , cmd_R89_ne996 , cmd_R89_ne997 , cmd_R89_ne297 : routeCommands;
	signal cmd_R30_Lc01 , cmd_R31_Lc01 , cmd_R32_Lc04 , cmd_R33_Lc04 : routeCommands;
	signal cmd_R2_D14 , cmd_R2_D15 , cmd_R3_D15 , cmd_R4_D18 , cmd_R4_D19 , cmd_R5_D19 , cmd_R6_D12 , cmd_R7_D12 , cmd_R8_D20 , cmd_R8_D21 , cmd_R9_D21 , cmd_R11_D04 , cmd_R11_Sw02 , cmd_R12_D15 , cmd_R13_D07 , cmd_R13_D16 , cmd_R14_D19 , cmd_R15_D21 , cmd_R16_D24 , cmd_R20_D01 , cmd_R21_Sw04 , cmd_R22_D14 , cmd_R26_D09 , cmd_R27_D23 , cmd_R28_D20 , cmd_R34_D05 , cmd_R35_D05 , cmd_R36_D05 , cmd_R37_D09 , cmd_R38_D09 , cmd_R39_D01 , cmd_R40_D01 , cmd_R41_D01 , cmd_R41_D03 , cmd_R42_D04 , cmd_R42_Sw02 , cmd_R43_D03 , cmd_R44_D03 , cmd_R45_D04 , cmd_R46_D04 , cmd_R47_D04 , cmd_R48_D07 , cmd_R49_D07 , cmd_R50_D07 , cmd_R51_D05 , cmd_R51_D08 , cmd_R52_D07 , cmd_R52_D16 , cmd_R53_D08 , cmd_R54_D08 , cmd_R55_D09 , cmd_R55_D10 , cmd_R56_D24 , cmd_R57_D10 , cmd_R58_D10 , cmd_R59_Sw02 , cmd_R60_D01 , cmd_R60_D03 , cmd_R60_Sw02 , cmd_R61_D14 , cmd_R62_D14 , cmd_R62_D15 , cmd_R63_D16 , cmd_R64_D05 , cmd_R64_D08 , cmd_R64_D16 , cmd_R65_D18 , cmd_R66_D18 , cmd_R67_D18 , cmd_R67_D19 , cmd_R68_D23 , cmd_R69_D23 , cmd_R69_D12 , cmd_R70_D23 , cmd_R70_D12 , cmd_R71_D23 , cmd_R71_D12 , cmd_R72_D12 , cmd_R73_D23 , cmd_R73_D12 , cmd_R74_D12 , cmd_R75_D20 , cmd_R75_D21 , cmd_R76_D20 , cmd_R77_D09 , cmd_R77_D10 , cmd_R77_D24 , cmd_R78_D24 , cmd_R79_Sw01 , cmd_R80_Sw01 , cmd_R81_Sw01 , cmd_R81_Sw05 , cmd_R82_Sw05 , cmd_R83_Sw05 , cmd_R84_Sw01 , cmd_R84_Sw05 , cmd_R85_Sw03 , cmd_R86_Sw03 , cmd_R87_Sw03 , cmd_R87_Sw04 , cmd_R88_Sw04 , cmd_R89_Sw03 , cmd_R89_Sw04 : routeCommands;
	signal cmd_R1_T02 , cmd_R2_T04 , cmd_R3_T04 , cmd_R4_T06 , cmd_R5_T06 , cmd_R6_T08 , cmd_R7_T08 , cmd_R8_T10 , cmd_R9_T10 , cmd_R10_T12 , cmd_R11_T14 , cmd_R12_T16 , cmd_R13_T18 , cmd_R14_T20 , cmd_R15_T22 , cmd_R16_T24 , cmd_R17_L29 , cmd_R18_L30 , cmd_R19_L31 , cmd_R20_J35 , cmd_R21_J36 , cmd_R22_J37 , cmd_R23_J38 , cmd_R24_J40 , cmd_R25_J43 , cmd_R26_J45 , cmd_R27_J46 , cmd_R28_J47 , cmd_R29_J48 , cmd_R30_X50 , cmd_R31_X51 , cmd_R32_X52 , cmd_R33_X53 , cmd_R34_C54 , cmd_R35_S55 , cmd_R36_S55 , cmd_R37_S59 , cmd_R38_S59 , cmd_R39_S64 , cmd_R40_S64 , cmd_R41_C67 , cmd_R42_B68 , cmd_R43_S69 , cmd_R44_S69 , cmd_R45_C70 , cmd_R46_S71 , cmd_R47_S71 , cmd_R48_C73 , cmd_R49_S74 , cmd_R50_S74 , cmd_R51_C76 , cmd_R52_B77 , cmd_R53_S78 , cmd_R54_S78 , cmd_R55_C79 , cmd_R56_B80 , cmd_R57_S81 , cmd_R58_S81 , cmd_R59_S84 , cmd_R60_S84 , cmd_R61_S86 , cmd_R62_S86 , cmd_R63_S93 , cmd_R64_S93 , cmd_R65_C94 , cmd_R66_S95 , cmd_R67_S95 , cmd_R68_S101 , cmd_R69_S101 , cmd_R70_S101 , cmd_R71_S104 , cmd_R72_S104 , cmd_R73_S107 , cmd_R74_S107 , cmd_R75_S110 , cmd_R76_S110 , cmd_R77_S117 , cmd_R78_S117 , cmd_R79_C119 , cmd_R80_S120 , cmd_R81_S120 , cmd_R82_C122 , cmd_R83_S123 , cmd_R84_S123 , cmd_R85_C125 , cmd_R86_S126 , cmd_R87_S126 , cmd_R88_S129 , cmd_R89_S129 : routeCommands;
begin
	levelCrossing_Lc01 : levelCrossing_0 port map(clock => clock, reset => reset, R30_command => cmd_R30_Lc01, R31_command => cmd_R31_Lc01, ocupation_ne98 => ocupation(20), ocupation_ne996 => ocupation(45), ocupation_ne99 => ocupation(21), indication => levelCrossings_i(0), command  => levelCrossings_o(0), lock_Lc01 => Lc01_locking, correspondence_Lc01 => state_Lc01);
	levelCrossing_Lc04 : levelCrossing_1 port map(clock => clock, reset => reset, R32_command => cmd_R32_Lc04, R33_command => cmd_R33_Lc04, ocupation_ne100 => ocupation(22), ocupation_ne992 => ocupation(41), ocupation_ne101 => ocupation(23), indication => levelCrossings_i(1), command  => levelCrossings_o(1), lock_Lc04 => Lc04_locking, correspondence_Lc04 => state_Lc04);
	singleSwitch_D01 : singleSwitch_0 port map(clock => clock, reset => reset, R20_command => cmd_R20_D01, R39_command => cmd_R39_D01, R40_command => cmd_R40_D01, R41_command => cmd_R41_D01, R60_command => cmd_R60_D01, indication => singleSwitches_i(0), command => singleSwitches_o(0), lock_D01 => D01_locking, correspondence_D01 => state_D01);
	singleSwitch_D08 : singleSwitch_1 port map(clock => clock, reset => reset, R51_command => cmd_R51_D08, R53_command => cmd_R53_D08, R54_command => cmd_R54_D08, R64_command => cmd_R64_D08, indication => singleSwitches_i(1), command => singleSwitches_o(1), lock_D08 => D08_locking, correspondence_D08 => state_D08);
	singleSwitch_D05 : singleSwitch_2 port map(clock => clock, reset => reset, R34_command => cmd_R34_D05, R35_command => cmd_R35_D05, R36_command => cmd_R36_D05, R51_command => cmd_R51_D05, R64_command => cmd_R64_D05, indication => singleSwitches_i(2), command => singleSwitches_o(2), lock_D05 => D05_locking, correspondence_D05 => state_D05);
	singleSwitch_D18 : singleSwitch_3 port map(clock => clock, reset => reset, R4_command => cmd_R4_D18, R65_command => cmd_R65_D18, R66_command => cmd_R66_D18, R67_command => cmd_R67_D18, indication => singleSwitches_i(3), command => singleSwitches_o(3), lock_D18 => D18_locking, correspondence_D18 => state_D18);
	singleSwitch_Sw01 : singleSwitch_4 port map(clock => clock, reset => reset, R79_command => cmd_R79_Sw01, R80_command => cmd_R80_Sw01, R81_command => cmd_R81_Sw01, R84_command => cmd_R84_Sw01, indication => singleSwitches_i(4), command => singleSwitches_o(4), lock_Sw01 => Sw01_locking, correspondence_Sw01 => state_Sw01);
	singleSwitch_D10 : singleSwitch_5 port map(clock => clock, reset => reset, R55_command => cmd_R55_D10, R57_command => cmd_R57_D10, R58_command => cmd_R58_D10, R77_command => cmd_R77_D10, indication => singleSwitches_i(5), command => singleSwitches_o(5), lock_D10 => D10_locking, correspondence_D10 => state_D10);
	singleSwitch_D09 : singleSwitch_6 port map(clock => clock, reset => reset, R26_command => cmd_R26_D09, R37_command => cmd_R37_D09, R38_command => cmd_R38_D09, R55_command => cmd_R55_D09, R77_command => cmd_R77_D09, indication => singleSwitches_i(6), command => singleSwitches_o(6), lock_D09 => D09_locking, correspondence_D09 => state_D09);
	singleSwitch_D20 : singleSwitch_7 port map(clock => clock, reset => reset, R8_command => cmd_R8_D20, R28_command => cmd_R28_D20, R75_command => cmd_R75_D20, R76_command => cmd_R76_D20, indication => singleSwitches_i(7), command => singleSwitches_o(7), lock_D20 => D20_locking, correspondence_D20 => state_D20);
	singleSwitch_D23 : singleSwitch_8 port map(clock => clock, reset => reset, R27_command => cmd_R27_D23, R68_command => cmd_R68_D23, R69_command => cmd_R69_D23, R70_command => cmd_R70_D23, R71_command => cmd_R71_D23, R73_command => cmd_R73_D23, indication => singleSwitches_i(8), command => singleSwitches_o(8), lock_D23 => D23_locking, correspondence_D23 => state_D23);
	singleSwitch_D03 : singleSwitch_9 port map(clock => clock, reset => reset, R41_command => cmd_R41_D03, R43_command => cmd_R43_D03, R44_command => cmd_R44_D03, R60_command => cmd_R60_D03, indication => singleSwitches_i(9), command => singleSwitches_o(9), lock_D03 => D03_locking, correspondence_D03 => state_D03);
	singleSwitch_D14 : singleSwitch_10 port map(clock => clock, reset => reset, R2_command => cmd_R2_D14, R22_command => cmd_R22_D14, R61_command => cmd_R61_D14, R62_command => cmd_R62_D14, indication => singleSwitches_i(10), command => singleSwitches_o(10), lock_D14 => D14_locking, correspondence_D14 => state_D14);
	singleSwitch_Sw04 : singleSwitch_11 port map(clock => clock, reset => reset, R21_command => cmd_R21_Sw04, R87_command => cmd_R87_Sw04, R88_command => cmd_R88_Sw04, R89_command => cmd_R89_Sw04, indication => singleSwitches_i(11), command => singleSwitches_o(11), lock_Sw04 => Sw04_locking, correspondence_Sw04 => state_Sw04);
	singleSwitch_D04 : singleSwitch_12 port map(clock => clock, reset => reset, R11_command => cmd_R11_D04, R42_command => cmd_R42_D04, R45_command => cmd_R45_D04, R46_command => cmd_R46_D04, R47_command => cmd_R47_D04, indication => singleSwitches_i(12), command => singleSwitches_o(12), lock_D04 => D04_locking, correspondence_D04 => state_D04);
	singleSwitch_Sw03 : singleSwitch_13 port map(clock => clock, reset => reset, R85_command => cmd_R85_Sw03, R86_command => cmd_R86_Sw03, R87_command => cmd_R87_Sw03, R89_command => cmd_R89_Sw03, indication => singleSwitches_i(13), command => singleSwitches_o(13), lock_Sw03 => Sw03_locking, correspondence_Sw03 => state_Sw03);
	singleSwitch_D15 : singleSwitch_14 port map(clock => clock, reset => reset, R2_command => cmd_R2_D15, R3_command => cmd_R3_D15, R12_command => cmd_R12_D15, R62_command => cmd_R62_D15, indication => singleSwitches_i(14), command => singleSwitches_o(14), lock_D15 => D15_locking, correspondence_D15 => state_D15);
	singleSwitch_Sw02 : singleSwitch_15 port map(clock => clock, reset => reset, R11_command => cmd_R11_Sw02, R42_command => cmd_R42_Sw02, R59_command => cmd_R59_Sw02, R60_command => cmd_R60_Sw02, indication => singleSwitches_i(15), command => singleSwitches_o(15), lock_Sw02 => Sw02_locking, correspondence_Sw02 => state_Sw02);
	singleSwitch_D07 : singleSwitch_16 port map(clock => clock, reset => reset, R13_command => cmd_R13_D07, R48_command => cmd_R48_D07, R49_command => cmd_R49_D07, R50_command => cmd_R50_D07, R52_command => cmd_R52_D07, indication => singleSwitches_i(16), command => singleSwitches_o(16), lock_D07 => D07_locking, correspondence_D07 => state_D07);
	singleSwitch_Sw05 : singleSwitch_17 port map(clock => clock, reset => reset, R81_command => cmd_R81_Sw05, R82_command => cmd_R82_Sw05, R83_command => cmd_R83_Sw05, R84_command => cmd_R84_Sw05, indication => singleSwitches_i(17), command => singleSwitches_o(17), lock_Sw05 => Sw05_locking, correspondence_Sw05 => state_Sw05);
	singleSwitch_D16 : singleSwitch_18 port map(clock => clock, reset => reset, R13_command => cmd_R13_D16, R52_command => cmd_R52_D16, R63_command => cmd_R63_D16, R64_command => cmd_R64_D16, indication => singleSwitches_i(18), command => singleSwitches_o(18), lock_D16 => D16_locking, correspondence_D16 => state_D16);
	singleSwitch_D19 : singleSwitch_19 port map(clock => clock, reset => reset, R4_command => cmd_R4_D19, R5_command => cmd_R5_D19, R14_command => cmd_R14_D19, R67_command => cmd_R67_D19, indication => singleSwitches_i(19), command => singleSwitches_o(19), lock_D19 => D19_locking, correspondence_D19 => state_D19);
	singleSwitch_D21 : singleSwitch_20 port map(clock => clock, reset => reset, R8_command => cmd_R8_D21, R9_command => cmd_R9_D21, R15_command => cmd_R15_D21, R75_command => cmd_R75_D21, indication => singleSwitches_i(20), command => singleSwitches_o(20), lock_D21 => D21_locking, correspondence_D21 => state_D21);
	singleSwitch_D24 : singleSwitch_21 port map(clock => clock, reset => reset, R16_command => cmd_R16_D24, R56_command => cmd_R56_D24, R77_command => cmd_R77_D24, R78_command => cmd_R78_D24, indication => singleSwitches_i(21), command => singleSwitches_o(21), lock_D24 => D24_locking, correspondence_D24 => state_D24);
	doubleSwitch_D12 : doubleSwitch_0 port map(clock => clock, reset => reset, R6_command => cmd_R6_D12, R7_command => cmd_R7_D12, R69_command => cmd_R69_D12, R70_command => cmd_R70_D12, R71_command => cmd_R71_D12, R72_command => cmd_R72_D12, R73_command => cmd_R73_D12, R74_command => cmd_R74_D12, indication => doubleSwitches_i, command => doubleSwitches_o, lock_D12 => D12_locking, correspondence_D12 => state_D12);
	railwaySignal_T01 : railwaySignal_0 port map(clock => clock, reset => reset, ocupation_ne991 => ocupation(0), indication.msb => signals_i.msb(0), indication.lsb => signals_i.lsb(0), command.msb => signals_o.msb(0), command.lsb => signals_o.lsb(0), lock_T01 => T01_locking, correspondence_T01 => state_T01);
	railwaySignal_T02 : railwaySignal_1 port map(clock => clock, reset => reset, R1_command => cmd_R1_T02, ocupation_ne991 => ocupation(0), ocupation_ne290 => ocupation(8), ocupation_ne288 => ocupation(7), correspondence_S64 => state_S64, correspondence_S69 => state_S69, correspondence_S86 => state_S86, D01_state => state_D01, indication.msb => signals_i.msb(1), indication.lsb => signals_i.lsb(1), command.msb => signals_o.msb(1), command.lsb => signals_o.lsb(1), lock_T02 => T02_locking, correspondence_T02 => state_T02);
	railwaySignal_S64 : railwaySignal_2 port map(clock => clock, reset => reset, R39_command => cmd_R39_S64, R40_command => cmd_R40_S64, ocupation_ne991 => ocupation(0), ocupation_ne288 => ocupation(7), ocupation_ne290 => ocupation(8), ocupation_ne110 => ocupation(26), ocupation_ne295 => ocupation(10), ocupation_ne111 => ocupation(27), ocupation_ne377 => ocupation(12), ocupation_ne292 => ocupation(9), correspondence_S69 => state_S69, correspondence_S86 => state_S86, correspondence_C70 => state_C70, correspondence_B68 => state_B68, correspondence_J36 => state_J36, correspondence_T03 => state_T03, D01_state => state_D01, D03_state => state_D03, D14_state => state_D14, D15_state => state_D15, indication.msb => signals_i.msb(2), indication.lsb => signals_i.lsb(2), command.msb => signals_o.msb(2), command.lsb => signals_o.lsb(2), lock_S64 => S64_locking, correspondence_S64 => state_S64);
	railwaySignal_S78 : railwaySignal_3 port map(clock => clock, reset => reset, R53_command => cmd_R53_S78, R54_command => cmd_R54_S78, ocupation_ne61 => ocupation(1), ocupation_ne404 => ocupation(15), ocupation_ne123 => ocupation(30), ocupation_ne400 => ocupation(14), ocupation_ne407 => ocupation(16), correspondence_C73 => state_C73, correspondence_B77 => state_B77, correspondence_S123 => state_S123, D08_state => state_D08, D07_state => state_D07, D16_state => state_D16, indication.msb => signals_i.msb(3), indication.lsb => signals_i.lsb(3), command.msb => signals_o.msb(3), command.lsb => signals_o.lsb(3), lock_S78 => S78_locking, correspondence_S78 => state_S78);
	railwaySignal_C54 : railwaySignal_4 port map(clock => clock, reset => reset, R34_command => cmd_R34_C54, ocupation_ne63 => ocupation(2), ocupation_ne99 => ocupation(21), ocupation_ne98 => ocupation(20), ocupation_ne996 => ocupation(45), correspondence_X51 => state_X51, correspondence_S129 => state_S129, D05_state => state_D05, Lc01_state => state_Lc01, indication.msb => signals_i.msb(4), indication.lsb => signals_i.lsb(4), command.msb => signals_o.msb(4), command.lsb => signals_o.lsb(4), lock_C54 => C54_locking, correspondence_C54 => state_C54);
	railwaySignal_S95 : railwaySignal_5 port map(clock => clock, reset => reset, R66_command => cmd_R66_S95, R67_command => cmd_R67_S95, ocupation_ne63 => ocupation(2), ocupation_ne65 => ocupation(3), ocupation_ne124 => ocupation(31), ocupation_ne421 => ocupation(17), ocupation_ne992 => ocupation(41), correspondence_C119 => state_C119, correspondence_T05 => state_T05, correspondence_J40 => state_J40, D18_state => state_D18, Sw01_state => state_Sw01, D19_state => state_D19, indication.msb => signals_i.msb(5), indication.lsb => signals_i.lsb(5), command.msb => signals_o.msb(5), command.lsb => signals_o.lsb(5), lock_S95 => S95_locking, correspondence_S95 => state_S95);
	railwaySignal_C94 : railwaySignal_6 port map(clock => clock, reset => reset, R65_command => cmd_R65_C94, ocupation_ne65 => ocupation(3), ocupation_ne63 => ocupation(2), ocupation_ne98 => ocupation(20), ocupation_ne99 => ocupation(21), correspondence_C54 => state_C54, correspondence_X51 => state_X51, D18_state => state_D18, D05_state => state_D05, indication.msb => signals_i.msb(6), indication.lsb => signals_i.lsb(6), command.msb => signals_o.msb(6), command.lsb => signals_o.lsb(6), lock_C94 => C94_locking, correspondence_C94 => state_C94);
	railwaySignal_C119 : railwaySignal_7 port map(clock => clock, reset => reset, R79_command => cmd_R79_C119, ocupation_ne65 => ocupation(3), ocupation_ne992 => ocupation(41), ocupation_ne100 => ocupation(22), correspondence_J40 => state_J40, correspondence_L31 => state_L31, Sw01_state => state_Sw01, indication.msb => signals_i.msb(7), indication.lsb => signals_i.lsb(7), command.msb => signals_o.msb(7), command.lsb => signals_o.lsb(7), lock_C119 => C119_locking, correspondence_C119 => state_C119);
	railwaySignal_S81 : railwaySignal_8 port map(clock => clock, reset => reset, R57_command => cmd_R57_S81, R58_command => cmd_R58_S81, ocupation_ne910 => ocupation(4), ocupation_ne130 => ocupation(35), ocupation_ne135 => ocupation(40), ocupation_ne114 => ocupation(6), ocupation_ne450 => ocupation(18), ocupation_ne129 => ocupation(34), ocupation_ne127 => ocupation(33), correspondence_S107 => state_S107, correspondence_B80 => state_B80, correspondence_L29 => state_L29, correspondence_T07 => state_T07, correspondence_S104 => state_S104, D10_state => state_D10, D23_state => state_D23, D12_state => state_D12, D24_state => state_D24, indication.msb => signals_i.msb(8), indication.lsb => signals_i.lsb(8), command.msb => signals_o.msb(8), command.lsb => signals_o.lsb(8), lock_S81 => S81_locking, correspondence_S81 => state_S81);
	railwaySignal_J45 : railwaySignal_9 port map(clock => clock, reset => reset, R26_command => cmd_R26_J45, ocupation_ne912 => ocupation(5), ocupation_ne101 => ocupation(23), ocupation_ne100 => ocupation(22), correspondence_J43 => state_J43, correspondence_X53 => state_X53, D09_state => state_D09, indication.msb => signals_i.msb(9), indication.lsb => signals_i.lsb(9), command.msb => signals_o.msb(9), command.lsb => signals_o.lsb(9), lock_J45 => J45_locking, correspondence_J45 => state_J45);
	railwaySignal_S110 : railwaySignal_10 port map(clock => clock, reset => reset, R75_command => cmd_R75_S110, R76_command => cmd_R76_S110, ocupation_ne912 => ocupation(5), ocupation_ne131 => ocupation(36), ocupation_ne465 => ocupation(19), ocupation_ne132 => ocupation(37), ocupation_ne114 => ocupation(6), correspondence_T09 => state_T09, correspondence_J46 => state_J46, correspondence_L29 => state_L29, D20_state => state_D20, D21_state => state_D21, D23_state => state_D23, indication.msb => signals_i.msb(10), indication.lsb => signals_i.lsb(10), command.msb => signals_o.msb(10), command.lsb => signals_o.lsb(10), lock_S110 => S110_locking, correspondence_S110 => state_S110);
	railwaySignal_L29 : railwaySignal_11 port map(clock => clock, reset => reset, R17_command => cmd_R17_L29, ocupation_ne114 => ocupation(6), ocupation_ne102 => ocupation(24), correspondence_J48 => state_J48, correspondence_T11 => state_T11, indication.msb => signals_i.msb(11), indication.lsb => signals_i.lsb(11), command.msb => signals_o.msb(11), command.lsb => signals_o.lsb(11), lock_L29 => L29_locking, correspondence_L29 => state_L29);
	railwaySignal_J48 : railwaySignal_12 port map(clock => clock, reset => reset, R29_command => cmd_R29_J48, ocupation_ne114 => ocupation(6), ocupation_ne102 => ocupation(24), correspondence_T11 => state_T11, indication.msb => signals_i.msb(12), indication.lsb => signals_i.lsb(12), command.msb => signals_o.msb(12), command.lsb => signals_o.lsb(12), lock_J48 => J48_locking, correspondence_J48 => state_J48);
	railwaySignal_S101 : railwaySignal_13 port map(clock => clock, reset => reset, R68_command => cmd_R68_S101, R69_command => cmd_R69_S101, R70_command => cmd_R70_S101, ocupation_ne114 => ocupation(6), ocupation_ne132 => ocupation(37), ocupation_ne129 => ocupation(34), ocupation_ne127 => ocupation(33), ocupation_ne130 => ocupation(35), ocupation_ne912 => ocupation(5), ocupation_ne910 => ocupation(4), ocupation_ne134 => ocupation(39), ocupation_ne135 => ocupation(40), ocupation_ne101 => ocupation(23), correspondence_J47 => state_J47, correspondence_S117 => state_S117, correspondence_C79 => state_C79, correspondence_J45 => state_J45, correspondence_J43 => state_J43, correspondence_T23 => state_T23, D23_state => state_D23, D20_state => state_D20, D12_state => state_D12, D09_state => state_D09, D10_state => state_D10, D24_state => state_D24, indication.msb => signals_i.msb(13), indication.lsb => signals_i.lsb(13), command.msb => signals_o.msb(13), command.lsb => signals_o.lsb(13), lock_S101 => S101_locking, correspondence_S101 => state_S101);
	railwaySignal_S69 : railwaySignal_14 port map(clock => clock, reset => reset, R43_command => cmd_R43_S69, R44_command => cmd_R44_S69, ocupation_ne288 => ocupation(7), ocupation_ne295 => ocupation(10), ocupation_ne110 => ocupation(26), ocupation_ne297 => ocupation(11), ocupation_ne384 => ocupation(13), correspondence_C70 => state_C70, correspondence_B68 => state_B68, correspondence_S126 => state_S126, D03_state => state_D03, D04_state => state_D04, Sw02_state => state_Sw02, indication.msb => signals_i.msb(14), indication.lsb => signals_i.lsb(14), command.msb => signals_o.msb(14), command.lsb => signals_o.lsb(14), lock_S69 => S69_locking, correspondence_S69 => state_S69);
	railwaySignal_J35 : railwaySignal_15 port map(clock => clock, reset => reset, R20_command => cmd_R20_J35, ocupation_ne290 => ocupation(8), ocupation_ne991 => ocupation(0), correspondence_T01 => state_T01, D01_state => state_D01, indication.msb => signals_i.msb(15), indication.lsb => signals_i.lsb(15), command.msb => signals_o.msb(15), command.lsb => signals_o.lsb(15), lock_J35 => J35_locking, correspondence_J35 => state_J35);
	railwaySignal_S86 : railwaySignal_16 port map(clock => clock, reset => reset, R61_command => cmd_R61_S86, R62_command => cmd_R62_S86, ocupation_ne290 => ocupation(8), ocupation_ne292 => ocupation(9), ocupation_ne111 => ocupation(27), ocupation_ne377 => ocupation(12), ocupation_ne996 => ocupation(45), correspondence_J36 => state_J36, correspondence_T03 => state_T03, correspondence_J38 => state_J38, D14_state => state_D14, Sw04_state => state_Sw04, D15_state => state_D15, indication.msb => signals_i.msb(16), indication.lsb => signals_i.lsb(16), command.msb => signals_o.msb(16), command.lsb => signals_o.lsb(16), lock_S86 => S86_locking, correspondence_S86 => state_S86);
	railwaySignal_J36 : railwaySignal_17 port map(clock => clock, reset => reset, R21_command => cmd_R21_J36, ocupation_ne292 => ocupation(9), ocupation_ne996 => ocupation(45), ocupation_ne98 => ocupation(20), correspondence_J38 => state_J38, correspondence_L30 => state_L30, Sw04_state => state_Sw04, indication.msb => signals_i.msb(17), indication.lsb => signals_i.lsb(17), command.msb => signals_o.msb(17), command.lsb => signals_o.lsb(17), lock_J36 => J36_locking, correspondence_J36 => state_J36);
	railwaySignal_J37 : railwaySignal_18 port map(clock => clock, reset => reset, R22_command => cmd_R22_J37, ocupation_ne292 => ocupation(9), ocupation_ne290 => ocupation(8), ocupation_ne991 => ocupation(0), correspondence_J35 => state_J35, correspondence_T01 => state_T01, D14_state => state_D14, D01_state => state_D01, indication.msb => signals_i.msb(18), indication.lsb => signals_i.lsb(18), command.msb => signals_o.msb(18), command.lsb => signals_o.lsb(18), lock_J37 => J37_locking, correspondence_J37 => state_J37);
	railwaySignal_C67 : railwaySignal_19 port map(clock => clock, reset => reset, R41_command => cmd_R41_C67, ocupation_ne295 => ocupation(10), ocupation_ne288 => ocupation(7), ocupation_ne991 => ocupation(0), correspondence_T01 => state_T01, D01_state => state_D01, D03_state => state_D03, indication.msb => signals_i.msb(19), indication.lsb => signals_i.lsb(19), command.msb => signals_o.msb(19), command.lsb => signals_o.lsb(19), lock_C67 => C67_locking, correspondence_C67 => state_C67);
	railwaySignal_C70 : railwaySignal_20 port map(clock => clock, reset => reset, R45_command => cmd_R45_C70, ocupation_ne295 => ocupation(10), ocupation_ne297 => ocupation(11), ocupation_ne996 => ocupation(45), ocupation_ne995 => ocupation(44), ocupation_ne997 => ocupation(46), correspondence_S126 => state_S126, correspondence_T27 => state_T27, correspondence_J38 => state_J38, D04_state => state_D04, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication.msb => signals_i.msb(20), indication.lsb => signals_i.lsb(20), command.msb => signals_o.msb(20), command.lsb => signals_o.lsb(20), lock_C70 => C70_locking, correspondence_C70 => state_C70);
	railwaySignal_S71 : railwaySignal_21 port map(clock => clock, reset => reset, R46_command => cmd_R46_S71, R47_command => cmd_R47_S71, ocupation_ne297 => ocupation(11), ocupation_ne295 => ocupation(10), ocupation_ne384 => ocupation(13), ocupation_ne991 => ocupation(0), ocupation_ne288 => ocupation(7), ocupation_ne110 => ocupation(26), ocupation_ne104 => ocupation(25), correspondence_C67 => state_C67, correspondence_S84 => state_S84, correspondence_T01 => state_T01, correspondence_T13 => state_T13, D04_state => state_D04, D01_state => state_D01, D03_state => state_D03, Sw02_state => state_Sw02, indication.msb => signals_i.msb(21), indication.lsb => signals_i.lsb(21), command.msb => signals_o.msb(21), command.lsb => signals_o.lsb(21), lock_S71 => S71_locking, correspondence_S71 => state_S71);
	railwaySignal_S126 : railwaySignal_22 port map(clock => clock, reset => reset, R86_command => cmd_R86_S126, R87_command => cmd_R87_S126, ocupation_ne297 => ocupation(11), ocupation_ne995 => ocupation(44), ocupation_ne997 => ocupation(46), ocupation_ne996 => ocupation(45), ocupation_ne98 => ocupation(20), correspondence_T27 => state_T27, correspondence_J38 => state_J38, correspondence_L30 => state_L30, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication.msb => signals_i.msb(22), indication.lsb => signals_i.lsb(22), command.msb => signals_o.msb(22), command.lsb => signals_o.lsb(22), lock_S126 => S126_locking, correspondence_S126 => state_S126);
	railwaySignal_T03 : railwaySignal_23 port map(clock => clock, reset => reset, ocupation_ne377 => ocupation(12), indication.msb => signals_i.msb(23), indication.lsb => signals_i.lsb(23), command.msb => signals_o.msb(23), command.lsb => signals_o.lsb(23), lock_T03 => T03_locking, correspondence_T03 => state_T03);
	railwaySignal_T04 : railwaySignal_24 port map(clock => clock, reset => reset, R2_command => cmd_R2_T04, R3_command => cmd_R3_T04, ocupation_ne377 => ocupation(12), ocupation_ne111 => ocupation(27), ocupation_ne290 => ocupation(8), ocupation_ne113 => ocupation(28), ocupation_ne991 => ocupation(0), correspondence_J35 => state_J35, correspondence_T15 => state_T15, correspondence_T01 => state_T01, D14_state => state_D14, D15_state => state_D15, D01_state => state_D01, indication.msb => signals_i.msb(24), indication.lsb => signals_i.lsb(24), command.msb => signals_o.msb(24), command.lsb => signals_o.lsb(24), lock_T04 => T04_locking, correspondence_T04 => state_T04);
	railwaySignal_S84 : railwaySignal_25 port map(clock => clock, reset => reset, R59_command => cmd_R59_S84, R60_command => cmd_R60_S84, ocupation_ne384 => ocupation(13), ocupation_ne104 => ocupation(25), ocupation_ne110 => ocupation(26), ocupation_ne288 => ocupation(7), ocupation_ne991 => ocupation(0), correspondence_T13 => state_T13, correspondence_T01 => state_T01, Sw02_state => state_Sw02, D01_state => state_D01, D03_state => state_D03, indication.msb => signals_i.msb(25), indication.lsb => signals_i.lsb(25), command.msb => signals_o.msb(25), command.lsb => signals_o.lsb(25), lock_S84 => S84_locking, correspondence_S84 => state_S84);
	railwaySignal_S74 : railwaySignal_26 port map(clock => clock, reset => reset, R49_command => cmd_R49_S74, R50_command => cmd_R50_S74, ocupation_ne400 => ocupation(14), ocupation_ne404 => ocupation(15), ocupation_ne407 => ocupation(16), ocupation_ne98 => ocupation(20), ocupation_ne99 => ocupation(21), ocupation_ne61 => ocupation(1), ocupation_ne123 => ocupation(30), ocupation_ne122 => ocupation(29), correspondence_C76 => state_C76, correspondence_S93 => state_S93, correspondence_X51 => state_X51, correspondence_T17 => state_T17, D07_state => state_D07, D05_state => state_D05, D08_state => state_D08, D16_state => state_D16, indication.msb => signals_i.msb(26), indication.lsb => signals_i.lsb(26), command.msb => signals_o.msb(26), command.lsb => signals_o.lsb(26), lock_S74 => S74_locking, correspondence_S74 => state_S74);
	railwaySignal_S123 : railwaySignal_27 port map(clock => clock, reset => reset, R83_command => cmd_R83_S123, R84_command => cmd_R84_S123, ocupation_ne400 => ocupation(14), ocupation_ne993 => ocupation(42), ocupation_ne994 => ocupation(43), ocupation_ne992 => ocupation(41), ocupation_ne100 => ocupation(22), correspondence_T25 => state_T25, correspondence_J40 => state_J40, correspondence_L31 => state_L31, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication.msb => signals_i.msb(27), indication.lsb => signals_i.lsb(27), command.msb => signals_o.msb(27), command.lsb => signals_o.lsb(27), lock_S123 => S123_locking, correspondence_S123 => state_S123);
	railwaySignal_C73 : railwaySignal_28 port map(clock => clock, reset => reset, R48_command => cmd_R48_C73, ocupation_ne404 => ocupation(15), ocupation_ne400 => ocupation(14), ocupation_ne992 => ocupation(41), ocupation_ne994 => ocupation(43), ocupation_ne993 => ocupation(42), correspondence_S123 => state_S123, correspondence_T25 => state_T25, correspondence_J40 => state_J40, D07_state => state_D07, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication.msb => signals_i.msb(28), indication.lsb => signals_i.lsb(28), command.msb => signals_o.msb(28), command.lsb => signals_o.lsb(28), lock_C73 => C73_locking, correspondence_C73 => state_C73);
	railwaySignal_C76 : railwaySignal_29 port map(clock => clock, reset => reset, R51_command => cmd_R51_C76, ocupation_ne404 => ocupation(15), ocupation_ne61 => ocupation(1), ocupation_ne99 => ocupation(21), ocupation_ne98 => ocupation(20), ocupation_ne996 => ocupation(45), correspondence_X51 => state_X51, correspondence_S129 => state_S129, D05_state => state_D05, D08_state => state_D08, Lc01_state => state_Lc01, indication.msb => signals_i.msb(29), indication.lsb => signals_i.lsb(29), command.msb => signals_o.msb(29), command.lsb => signals_o.lsb(29), lock_C76 => C76_locking, correspondence_C76 => state_C76);
	railwaySignal_S93 : railwaySignal_30 port map(clock => clock, reset => reset, R63_command => cmd_R63_S93, R64_command => cmd_R64_S93, ocupation_ne407 => ocupation(16), ocupation_ne122 => ocupation(29), ocupation_ne123 => ocupation(30), ocupation_ne61 => ocupation(1), ocupation_ne99 => ocupation(21), ocupation_ne98 => ocupation(20), ocupation_ne996 => ocupation(45), correspondence_T17 => state_T17, correspondence_X51 => state_X51, correspondence_S129 => state_S129, D16_state => state_D16, D05_state => state_D05, D08_state => state_D08, Lc01_state => state_Lc01, indication.msb => signals_i.msb(30), indication.lsb => signals_i.lsb(30), command.msb => signals_o.msb(30), command.lsb => signals_o.lsb(30), lock_S93 => S93_locking, correspondence_S93 => state_S93);
	railwaySignal_T05 : railwaySignal_31 port map(clock => clock, reset => reset, ocupation_ne421 => ocupation(17), indication.msb => signals_i.msb(31), indication.lsb => signals_i.lsb(31), command.msb => signals_o.msb(31), command.lsb => signals_o.lsb(31), lock_T05 => T05_locking, correspondence_T05 => state_T05);
	railwaySignal_T06 : railwaySignal_32 port map(clock => clock, reset => reset, R4_command => cmd_R4_T06, R5_command => cmd_R5_T06, ocupation_ne421 => ocupation(17), ocupation_ne124 => ocupation(31), ocupation_ne63 => ocupation(2), ocupation_ne126 => ocupation(32), ocupation_ne98 => ocupation(20), ocupation_ne99 => ocupation(21), correspondence_C54 => state_C54, correspondence_T19 => state_T19, correspondence_X51 => state_X51, D18_state => state_D18, D19_state => state_D19, D05_state => state_D05, indication.msb => signals_i.msb(32), indication.lsb => signals_i.lsb(32), command.msb => signals_o.msb(32), command.lsb => signals_o.lsb(32), lock_T06 => T06_locking, correspondence_T06 => state_T06);
	railwaySignal_T07 : railwaySignal_33 port map(clock => clock, reset => reset, ocupation_ne450 => ocupation(18), indication.msb => signals_i.msb(33), indication.lsb => signals_i.lsb(33), command.msb => signals_o.msb(33), command.lsb => signals_o.lsb(33), lock_T07 => T07_locking, correspondence_T07 => state_T07);
	railwaySignal_T08 : railwaySignal_34 port map(clock => clock, reset => reset, R6_command => cmd_R6_T08, R7_command => cmd_R7_T08, ocupation_ne450 => ocupation(18), ocupation_ne127 => ocupation(33), ocupation_ne130 => ocupation(35), ocupation_ne910 => ocupation(4), ocupation_ne134 => ocupation(39), ocupation_ne135 => ocupation(40), ocupation_ne101 => ocupation(23), correspondence_S117 => state_S117, correspondence_C79 => state_C79, correspondence_J43 => state_J43, correspondence_T23 => state_T23, D12_state => state_D12, D09_state => state_D09, D10_state => state_D10, D24_state => state_D24, indication.msb => signals_i.msb(34), indication.lsb => signals_i.lsb(34), command.msb => signals_o.msb(34), command.lsb => signals_o.lsb(34), lock_T08 => T08_locking, correspondence_T08 => state_T08);
	railwaySignal_T09 : railwaySignal_35 port map(clock => clock, reset => reset, ocupation_ne465 => ocupation(19), indication.msb => signals_i.msb(35), indication.lsb => signals_i.lsb(35), command.msb => signals_o.msb(35), command.lsb => signals_o.lsb(35), lock_T09 => T09_locking, correspondence_T09 => state_T09);
	railwaySignal_T10 : railwaySignal_36 port map(clock => clock, reset => reset, R8_command => cmd_R8_T10, R9_command => cmd_R9_T10, ocupation_ne465 => ocupation(19), ocupation_ne131 => ocupation(36), ocupation_ne912 => ocupation(5), ocupation_ne133 => ocupation(38), ocupation_ne101 => ocupation(23), correspondence_J45 => state_J45, correspondence_T21 => state_T21, correspondence_J43 => state_J43, D20_state => state_D20, D21_state => state_D21, D09_state => state_D09, indication.msb => signals_i.msb(36), indication.lsb => signals_i.lsb(36), command.msb => signals_o.msb(36), command.lsb => signals_o.lsb(36), lock_T10 => T10_locking, correspondence_T10 => state_T10);
	railwaySignal_L30 : railwaySignal_37 port map(clock => clock, reset => reset, R18_command => cmd_R18_L30, ocupation_ne98 => ocupation(20), ocupation_ne99 => ocupation(21), correspondence_X50 => state_X50, correspondence_S55 => state_S55, indication.msb => signals_i.msb(37), indication.lsb => signals_i.lsb(37), command.msb => signals_o.msb(37), command.lsb => signals_o.lsb(37), lock_L30 => L30_locking, correspondence_L30 => state_L30);
	railwaySignal_X50 : railwaySignal_38 port map(clock => clock, reset => reset, R30_command => cmd_R30_X50, ocupation_ne98 => ocupation(20), ocupation_ne99 => ocupation(21), ocupation_ne61 => ocupation(1), ocupation_ne63 => ocupation(2), correspondence_S55 => state_S55, correspondence_S78 => state_S78, correspondence_S95 => state_S95, D05_state => state_D05, Lc01_state => state_Lc01, indication.msb => signals_i.msb(38), indication.lsb => signals_i.lsb(38), command.msb => signals_o.msb(38), command.lsb => signals_o.lsb(38), lock_X50 => X50_locking, correspondence_X50 => state_X50);
	railwaySignal_X51 : railwaySignal_39 port map(clock => clock, reset => reset, R31_command => cmd_R31_X51, ocupation_ne98 => ocupation(20), ocupation_ne996 => ocupation(45), ocupation_ne297 => ocupation(11), ocupation_ne292 => ocupation(9), ocupation_ne997 => ocupation(46), correspondence_S129 => state_S129, correspondence_J37 => state_J37, correspondence_S71 => state_S71, Sw04_state => state_Sw04, Sw03_state => state_Sw03, Lc01_state => state_Lc01, indication.msb => signals_i.msb(39), indication.lsb => signals_i.lsb(39), command.msb => signals_o.msb(39), command.lsb => signals_o.lsb(39), lock_X51 => X51_locking, correspondence_X51 => state_X51);
	railwaySignal_S55 : railwaySignal_40 port map(clock => clock, reset => reset, R35_command => cmd_R35_S55, R36_command => cmd_R36_S55, ocupation_ne99 => ocupation(21), ocupation_ne61 => ocupation(1), ocupation_ne63 => ocupation(2), ocupation_ne123 => ocupation(30), ocupation_ne404 => ocupation(15), ocupation_ne421 => ocupation(17), ocupation_ne65 => ocupation(3), ocupation_ne124 => ocupation(31), correspondence_S78 => state_S78, correspondence_S95 => state_S95, correspondence_C73 => state_C73, correspondence_B77 => state_B77, correspondence_C119 => state_C119, correspondence_T05 => state_T05, D05_state => state_D05, D08_state => state_D08, D18_state => state_D18, D19_state => state_D19, indication.msb => signals_i.msb(40), indication.lsb => signals_i.lsb(40), command.msb => signals_o.msb(40), command.lsb => signals_o.lsb(40), lock_S55 => S55_locking, correspondence_S55 => state_S55);
	railwaySignal_L31 : railwaySignal_41 port map(clock => clock, reset => reset, R19_command => cmd_R19_L31, ocupation_ne100 => ocupation(22), ocupation_ne101 => ocupation(23), correspondence_X52 => state_X52, correspondence_S59 => state_S59, indication.msb => signals_i.msb(41), indication.lsb => signals_i.lsb(41), command.msb => signals_o.msb(41), command.lsb => signals_o.lsb(41), lock_L31 => L31_locking, correspondence_L31 => state_L31);
	railwaySignal_X52 : railwaySignal_42 port map(clock => clock, reset => reset, R32_command => cmd_R32_X52, ocupation_ne100 => ocupation(22), ocupation_ne101 => ocupation(23), ocupation_ne910 => ocupation(4), ocupation_ne912 => ocupation(5), correspondence_S59 => state_S59, correspondence_S110 => state_S110, correspondence_S81 => state_S81, D09_state => state_D09, Lc04_state => state_Lc04, indication.msb => signals_i.msb(42), indication.lsb => signals_i.lsb(42), command.msb => signals_o.msb(42), command.lsb => signals_o.lsb(42), lock_X52 => X52_locking, correspondence_X52 => state_X52);
	railwaySignal_X53 : railwaySignal_43 port map(clock => clock, reset => reset, R33_command => cmd_R33_X53, ocupation_ne100 => ocupation(22), ocupation_ne992 => ocupation(41), ocupation_ne65 => ocupation(3), ocupation_ne994 => ocupation(43), ocupation_ne400 => ocupation(14), correspondence_S120 => state_S120, correspondence_C94 => state_C94, correspondence_S74 => state_S74, Sw01_state => state_Sw01, Sw05_state => state_Sw05, Lc04_state => state_Lc04, indication.msb => signals_i.msb(43), indication.lsb => signals_i.lsb(43), command.msb => signals_o.msb(43), command.lsb => signals_o.lsb(43), lock_X53 => X53_locking, correspondence_X53 => state_X53);
	railwaySignal_J43 : railwaySignal_44 port map(clock => clock, reset => reset, R25_command => cmd_R25_J43, ocupation_ne101 => ocupation(23), ocupation_ne100 => ocupation(22), ocupation_ne992 => ocupation(41), correspondence_X53 => state_X53, correspondence_S120 => state_S120, indication.msb => signals_i.msb(44), indication.lsb => signals_i.lsb(44), command.msb => signals_o.msb(44), command.lsb => signals_o.lsb(44), lock_J43 => J43_locking, correspondence_J43 => state_J43);
	railwaySignal_S59 : railwaySignal_45 port map(clock => clock, reset => reset, R37_command => cmd_R37_S59, R38_command => cmd_R38_S59, ocupation_ne101 => ocupation(23), ocupation_ne912 => ocupation(5), ocupation_ne910 => ocupation(4), ocupation_ne132 => ocupation(37), ocupation_ne465 => ocupation(19), ocupation_ne131 => ocupation(36), ocupation_ne130 => ocupation(35), ocupation_ne135 => ocupation(40), correspondence_S110 => state_S110, correspondence_S81 => state_S81, correspondence_T09 => state_T09, correspondence_J46 => state_J46, correspondence_S107 => state_S107, correspondence_B80 => state_B80, D09_state => state_D09, D20_state => state_D20, D21_state => state_D21, D10_state => state_D10, indication.msb => signals_i.msb(45), indication.lsb => signals_i.lsb(45), command.msb => signals_o.msb(45), command.lsb => signals_o.lsb(45), lock_S59 => S59_locking, correspondence_S59 => state_S59);
	railwaySignal_T11 : railwaySignal_46 port map(clock => clock, reset => reset, ocupation_ne102 => ocupation(24), indication.msb => signals_i.msb(46), indication.lsb => signals_i.lsb(46), command.msb => signals_o.msb(46), command.lsb => signals_o.lsb(46), lock_T11 => T11_locking, correspondence_T11 => state_T11);
	railwaySignal_T12 : railwaySignal_47 port map(clock => clock, reset => reset, R10_command => cmd_R10_T12, ocupation_ne102 => ocupation(24), ocupation_ne114 => ocupation(6), ocupation_ne132 => ocupation(37), ocupation_ne130 => ocupation(35), ocupation_ne127 => ocupation(33), ocupation_ne129 => ocupation(34), correspondence_S101 => state_S101, correspondence_J47 => state_J47, correspondence_S117 => state_S117, correspondence_C79 => state_C79, D23_state => state_D23, D12_state => state_D12, indication.msb => signals_i.msb(47), indication.lsb => signals_i.lsb(47), command.msb => signals_o.msb(47), command.lsb => signals_o.lsb(47), lock_T12 => T12_locking, correspondence_T12 => state_T12);
	railwaySignal_T13 : railwaySignal_48 port map(clock => clock, reset => reset, ocupation_ne104 => ocupation(25), indication.msb => signals_i.msb(48), indication.lsb => signals_i.lsb(48), command.msb => signals_o.msb(48), command.lsb => signals_o.lsb(48), lock_T13 => T13_locking, correspondence_T13 => state_T13);
	railwaySignal_T14 : railwaySignal_49 port map(clock => clock, reset => reset, R11_command => cmd_R11_T14, ocupation_ne104 => ocupation(25), ocupation_ne384 => ocupation(13), ocupation_ne297 => ocupation(11), ocupation_ne996 => ocupation(45), ocupation_ne995 => ocupation(44), ocupation_ne997 => ocupation(46), correspondence_S126 => state_S126, correspondence_T27 => state_T27, correspondence_J38 => state_J38, D04_state => state_D04, Sw02_state => state_Sw02, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication.msb => signals_i.msb(49), indication.lsb => signals_i.lsb(49), command.msb => signals_o.msb(49), command.lsb => signals_o.lsb(49), lock_T14 => T14_locking, correspondence_T14 => state_T14);
	railwaySignal_B68 : railwaySignal_50 port map(clock => clock, reset => reset, R42_command => cmd_R42_B68, ocupation_ne110 => ocupation(26), ocupation_ne384 => ocupation(13), ocupation_ne297 => ocupation(11), ocupation_ne996 => ocupation(45), ocupation_ne995 => ocupation(44), ocupation_ne997 => ocupation(46), correspondence_S126 => state_S126, correspondence_T27 => state_T27, correspondence_J38 => state_J38, D04_state => state_D04, Sw02_state => state_Sw02, Sw03_state => state_Sw03, Sw04_state => state_Sw04, indication.msb => signals_i.msb(50), indication.lsb => signals_i.lsb(50), command.msb => signals_o.msb(50), command.lsb => signals_o.lsb(50), lock_B68 => B68_locking, correspondence_B68 => state_B68);
	railwaySignal_T15 : railwaySignal_51 port map(clock => clock, reset => reset, ocupation_ne113 => ocupation(28), indication.msb => signals_i.msb(51), indication.lsb => signals_i.lsb(51), command.msb => signals_o.msb(51), command.lsb => signals_o.lsb(51), lock_T15 => T15_locking, correspondence_T15 => state_T15);
	railwaySignal_T16 : railwaySignal_52 port map(clock => clock, reset => reset, R12_command => cmd_R12_T16, ocupation_ne113 => ocupation(28), ocupation_ne377 => ocupation(12), correspondence_T03 => state_T03, D15_state => state_D15, indication.msb => signals_i.msb(52), indication.lsb => signals_i.lsb(52), command.msb => signals_o.msb(52), command.lsb => signals_o.lsb(52), lock_T16 => T16_locking, correspondence_T16 => state_T16);
	railwaySignal_T17 : railwaySignal_53 port map(clock => clock, reset => reset, ocupation_ne122 => ocupation(29), indication.msb => signals_i.msb(53), indication.lsb => signals_i.lsb(53), command.msb => signals_o.msb(53), command.lsb => signals_o.lsb(53), lock_T17 => T17_locking, correspondence_T17 => state_T17);
	railwaySignal_T18 : railwaySignal_54 port map(clock => clock, reset => reset, R13_command => cmd_R13_T18, ocupation_ne122 => ocupation(29), ocupation_ne407 => ocupation(16), ocupation_ne400 => ocupation(14), ocupation_ne992 => ocupation(41), ocupation_ne994 => ocupation(43), ocupation_ne993 => ocupation(42), correspondence_S123 => state_S123, correspondence_T25 => state_T25, correspondence_J40 => state_J40, D07_state => state_D07, D16_state => state_D16, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication.msb => signals_i.msb(54), indication.lsb => signals_i.lsb(54), command.msb => signals_o.msb(54), command.lsb => signals_o.lsb(54), lock_T18 => T18_locking, correspondence_T18 => state_T18);
	railwaySignal_B77 : railwaySignal_55 port map(clock => clock, reset => reset, R52_command => cmd_R52_B77, ocupation_ne123 => ocupation(30), ocupation_ne407 => ocupation(16), ocupation_ne400 => ocupation(14), ocupation_ne992 => ocupation(41), ocupation_ne994 => ocupation(43), ocupation_ne993 => ocupation(42), correspondence_S123 => state_S123, correspondence_T25 => state_T25, correspondence_J40 => state_J40, D07_state => state_D07, D16_state => state_D16, Sw05_state => state_Sw05, Sw01_state => state_Sw01, indication.msb => signals_i.msb(55), indication.lsb => signals_i.lsb(55), command.msb => signals_o.msb(55), command.lsb => signals_o.lsb(55), lock_B77 => B77_locking, correspondence_B77 => state_B77);
	railwaySignal_T19 : railwaySignal_56 port map(clock => clock, reset => reset, ocupation_ne126 => ocupation(32), indication.msb => signals_i.msb(56), indication.lsb => signals_i.lsb(56), command.msb => signals_o.msb(56), command.lsb => signals_o.lsb(56), lock_T19 => T19_locking, correspondence_T19 => state_T19);
	railwaySignal_T20 : railwaySignal_57 port map(clock => clock, reset => reset, R14_command => cmd_R14_T20, ocupation_ne126 => ocupation(32), ocupation_ne421 => ocupation(17), correspondence_T05 => state_T05, D19_state => state_D19, indication.msb => signals_i.msb(57), indication.lsb => signals_i.lsb(57), command.msb => signals_o.msb(57), command.lsb => signals_o.lsb(57), lock_T20 => T20_locking, correspondence_T20 => state_T20);
	railwaySignal_S104 : railwaySignal_58 port map(clock => clock, reset => reset, R71_command => cmd_R71_S104, R72_command => cmd_R72_S104, ocupation_ne127 => ocupation(33), ocupation_ne129 => ocupation(34), ocupation_ne114 => ocupation(6), ocupation_ne450 => ocupation(18), correspondence_L29 => state_L29, correspondence_T07 => state_T07, correspondence_J48 => state_J48, D23_state => state_D23, D12_state => state_D12, indication.msb => signals_i.msb(58), indication.lsb => signals_i.lsb(58), command.msb => signals_o.msb(58), command.lsb => signals_o.lsb(58), lock_S104 => S104_locking, correspondence_S104 => state_S104);
	railwaySignal_S117 : railwaySignal_59 port map(clock => clock, reset => reset, R77_command => cmd_R77_S117, R78_command => cmd_R78_S117, ocupation_ne127 => ocupation(33), ocupation_ne135 => ocupation(40), ocupation_ne910 => ocupation(4), ocupation_ne101 => ocupation(23), ocupation_ne134 => ocupation(39), ocupation_ne100 => ocupation(22), correspondence_J43 => state_J43, correspondence_T23 => state_T23, correspondence_X53 => state_X53, D09_state => state_D09, D10_state => state_D10, D24_state => state_D24, indication.msb => signals_i.msb(59), indication.lsb => signals_i.lsb(59), command.msb => signals_o.msb(59), command.lsb => signals_o.lsb(59), lock_S117 => S117_locking, correspondence_S117 => state_S117);
	railwaySignal_C79 : railwaySignal_60 port map(clock => clock, reset => reset, R55_command => cmd_R55_C79, ocupation_ne130 => ocupation(35), ocupation_ne910 => ocupation(4), ocupation_ne101 => ocupation(23), ocupation_ne100 => ocupation(22), correspondence_J43 => state_J43, correspondence_X53 => state_X53, D09_state => state_D09, D10_state => state_D10, indication.msb => signals_i.msb(60), indication.lsb => signals_i.lsb(60), command.msb => signals_o.msb(60), command.lsb => signals_o.lsb(60), lock_C79 => C79_locking, correspondence_C79 => state_C79);
	railwaySignal_S107 : railwaySignal_61 port map(clock => clock, reset => reset, R73_command => cmd_R73_S107, R74_command => cmd_R74_S107, ocupation_ne130 => ocupation(35), ocupation_ne129 => ocupation(34), ocupation_ne114 => ocupation(6), ocupation_ne450 => ocupation(18), correspondence_L29 => state_L29, correspondence_T07 => state_T07, correspondence_J48 => state_J48, D23_state => state_D23, D12_state => state_D12, indication.msb => signals_i.msb(61), indication.lsb => signals_i.lsb(61), command.msb => signals_o.msb(61), command.lsb => signals_o.lsb(61), lock_S107 => S107_locking, correspondence_S107 => state_S107);
	railwaySignal_J46 : railwaySignal_62 port map(clock => clock, reset => reset, R27_command => cmd_R27_J46, ocupation_ne132 => ocupation(37), ocupation_ne114 => ocupation(6), correspondence_L29 => state_L29, correspondence_J48 => state_J48, D23_state => state_D23, indication.msb => signals_i.msb(62), indication.lsb => signals_i.lsb(62), command.msb => signals_o.msb(62), command.lsb => signals_o.lsb(62), lock_J46 => J46_locking, correspondence_J46 => state_J46);
	railwaySignal_J47 : railwaySignal_63 port map(clock => clock, reset => reset, R28_command => cmd_R28_J47, ocupation_ne132 => ocupation(37), ocupation_ne912 => ocupation(5), ocupation_ne101 => ocupation(23), correspondence_J45 => state_J45, correspondence_J43 => state_J43, D20_state => state_D20, D09_state => state_D09, indication.msb => signals_i.msb(63), indication.lsb => signals_i.lsb(63), command.msb => signals_o.msb(63), command.lsb => signals_o.lsb(63), lock_J47 => J47_locking, correspondence_J47 => state_J47);
	railwaySignal_T21 : railwaySignal_64 port map(clock => clock, reset => reset, ocupation_ne133 => ocupation(38), indication.msb => signals_i.msb(64), indication.lsb => signals_i.lsb(64), command.msb => signals_o.msb(64), command.lsb => signals_o.lsb(64), lock_T21 => T21_locking, correspondence_T21 => state_T21);
	railwaySignal_T22 : railwaySignal_65 port map(clock => clock, reset => reset, R15_command => cmd_R15_T22, ocupation_ne133 => ocupation(38), ocupation_ne465 => ocupation(19), correspondence_T09 => state_T09, D21_state => state_D21, indication.msb => signals_i.msb(65), indication.lsb => signals_i.lsb(65), command.msb => signals_o.msb(65), command.lsb => signals_o.lsb(65), lock_T22 => T22_locking, correspondence_T22 => state_T22);
	railwaySignal_T23 : railwaySignal_66 port map(clock => clock, reset => reset, ocupation_ne134 => ocupation(39), indication.msb => signals_i.msb(66), indication.lsb => signals_i.lsb(66), command.msb => signals_o.msb(66), command.lsb => signals_o.lsb(66), lock_T23 => T23_locking, correspondence_T23 => state_T23);
	railwaySignal_T24 : railwaySignal_67 port map(clock => clock, reset => reset, R16_command => cmd_R16_T24, ocupation_ne134 => ocupation(39), ocupation_ne127 => ocupation(33), ocupation_ne114 => ocupation(6), ocupation_ne450 => ocupation(18), ocupation_ne129 => ocupation(34), correspondence_S104 => state_S104, correspondence_L29 => state_L29, correspondence_T07 => state_T07, D24_state => state_D24, D23_state => state_D23, D12_state => state_D12, indication.msb => signals_i.msb(67), indication.lsb => signals_i.lsb(67), command.msb => signals_o.msb(67), command.lsb => signals_o.lsb(67), lock_T24 => T24_locking, correspondence_T24 => state_T24);
	railwaySignal_B80 : railwaySignal_68 port map(clock => clock, reset => reset, R56_command => cmd_R56_B80, ocupation_ne135 => ocupation(40), ocupation_ne127 => ocupation(33), ocupation_ne114 => ocupation(6), ocupation_ne450 => ocupation(18), ocupation_ne129 => ocupation(34), correspondence_S104 => state_S104, correspondence_L29 => state_L29, correspondence_T07 => state_T07, D24_state => state_D24, D23_state => state_D23, D12_state => state_D12, indication.msb => signals_i.msb(68), indication.lsb => signals_i.lsb(68), command.msb => signals_o.msb(68), command.lsb => signals_o.lsb(68), lock_B80 => B80_locking, correspondence_B80 => state_B80);
	railwaySignal_J40 : railwaySignal_69 port map(clock => clock, reset => reset, R24_command => cmd_R24_J40, ocupation_ne992 => ocupation(41), ocupation_ne100 => ocupation(22), correspondence_L31 => state_L31, correspondence_X52 => state_X52, indication.msb => signals_i.msb(69), indication.lsb => signals_i.lsb(69), command.msb => signals_o.msb(69), command.lsb => signals_o.lsb(69), lock_J40 => J40_locking, correspondence_J40 => state_J40);
	railwaySignal_S120 : railwaySignal_70 port map(clock => clock, reset => reset, R80_command => cmd_R80_S120, R81_command => cmd_R81_S120, ocupation_ne992 => ocupation(41), ocupation_ne65 => ocupation(3), ocupation_ne994 => ocupation(43), ocupation_ne400 => ocupation(14), ocupation_ne63 => ocupation(2), ocupation_ne407 => ocupation(16), ocupation_ne404 => ocupation(15), correspondence_C94 => state_C94, correspondence_S74 => state_S74, correspondence_C54 => state_C54, correspondence_C76 => state_C76, correspondence_S93 => state_S93, Sw01_state => state_Sw01, D18_state => state_D18, Sw05_state => state_Sw05, D07_state => state_D07, indication.msb => signals_i.msb(70), indication.lsb => signals_i.lsb(70), command.msb => signals_o.msb(70), command.lsb => signals_o.lsb(70), lock_S120 => S120_locking, correspondence_S120 => state_S120);
	railwaySignal_T25 : railwaySignal_71 port map(clock => clock, reset => reset, ocupation_ne993 => ocupation(42), indication.msb => signals_i.msb(71), indication.lsb => signals_i.lsb(71), command.msb => signals_o.msb(71), command.lsb => signals_o.lsb(71), lock_T25 => T25_locking, correspondence_T25 => state_T25);
	railwaySignal_C122 : railwaySignal_72 port map(clock => clock, reset => reset, R82_command => cmd_R82_C122, ocupation_ne993 => ocupation(42), ocupation_ne400 => ocupation(14), ocupation_ne407 => ocupation(16), ocupation_ne404 => ocupation(15), correspondence_S74 => state_S74, correspondence_C76 => state_C76, correspondence_S93 => state_S93, Sw05_state => state_Sw05, D07_state => state_D07, indication.msb => signals_i.msb(72), indication.lsb => signals_i.lsb(72), command.msb => signals_o.msb(72), command.lsb => signals_o.lsb(72), lock_C122 => C122_locking, correspondence_C122 => state_C122);
	railwaySignal_T27 : railwaySignal_73 port map(clock => clock, reset => reset, ocupation_ne995 => ocupation(44), indication.msb => signals_i.msb(73), indication.lsb => signals_i.lsb(73), command.msb => signals_o.msb(73), command.lsb => signals_o.lsb(73), lock_T27 => T27_locking, correspondence_T27 => state_T27);
	railwaySignal_C125 : railwaySignal_74 port map(clock => clock, reset => reset, R85_command => cmd_R85_C125, ocupation_ne995 => ocupation(44), ocupation_ne297 => ocupation(11), ocupation_ne384 => ocupation(13), ocupation_ne295 => ocupation(10), correspondence_S71 => state_S71, correspondence_C67 => state_C67, correspondence_S84 => state_S84, Sw03_state => state_Sw03, D04_state => state_D04, indication.msb => signals_i.msb(74), indication.lsb => signals_i.lsb(74), command.msb => signals_o.msb(74), command.lsb => signals_o.lsb(74), lock_C125 => C125_locking, correspondence_C125 => state_C125);
	railwaySignal_J38 : railwaySignal_75 port map(clock => clock, reset => reset, R23_command => cmd_R23_J38, ocupation_ne996 => ocupation(45), ocupation_ne98 => ocupation(20), correspondence_L30 => state_L30, correspondence_X50 => state_X50, indication.msb => signals_i.msb(75), indication.lsb => signals_i.lsb(75), command.msb => signals_o.msb(75), command.lsb => signals_o.lsb(75), lock_J38 => J38_locking, correspondence_J38 => state_J38);
	railwaySignal_S129 : railwaySignal_76 port map(clock => clock, reset => reset, R88_command => cmd_R88_S129, R89_command => cmd_R89_S129, ocupation_ne996 => ocupation(45), ocupation_ne292 => ocupation(9), ocupation_ne997 => ocupation(46), ocupation_ne297 => ocupation(11), ocupation_ne290 => ocupation(8), ocupation_ne384 => ocupation(13), ocupation_ne295 => ocupation(10), correspondence_J37 => state_J37, correspondence_S71 => state_S71, correspondence_J35 => state_J35, correspondence_C67 => state_C67, correspondence_S84 => state_S84, Sw04_state => state_Sw04, D14_state => state_D14, Sw03_state => state_Sw03, D04_state => state_D04, indication.msb => signals_i.msb(76), indication.lsb => signals_i.lsb(76), command.msb => signals_o.msb(76), command.lsb => signals_o.lsb(76), lock_S129 => S129_locking, correspondence_S129 => state_S129);
	node_ne991 : node_0 port map(clock => clock, ocupation => ocupation(0), reset => reset, R1_command => cmd_R1_ne991, R20_command => cmd_R20_ne991, R39_command => cmd_R39_ne991, R40_command => cmd_R40_ne991, R41_command => cmd_R41_ne991, R60_command => cmd_R60_ne991, state => state_ne991, locking => ne991_locking);
	node_ne61 : node_1 port map(clock => clock, ocupation => ocupation(1), reset => reset, R35_command => cmd_R35_ne61, R51_command => cmd_R51_ne61, R53_command => cmd_R53_ne61, R54_command => cmd_R54_ne61, R64_command => cmd_R64_ne61, state => state_ne61, locking => ne61_locking);
	node_ne63 : node_2 port map(clock => clock, ocupation => ocupation(2), reset => reset, R4_command => cmd_R4_ne63, R34_command => cmd_R34_ne63, R36_command => cmd_R36_ne63, R65_command => cmd_R65_ne63, R66_command => cmd_R66_ne63, R67_command => cmd_R67_ne63, state => state_ne63, locking => ne63_locking);
	node_ne65 : node_3 port map(clock => clock, ocupation => ocupation(3), reset => reset, R65_command => cmd_R65_ne65, R66_command => cmd_R66_ne65, R79_command => cmd_R79_ne65, R80_command => cmd_R80_ne65, state => state_ne65, locking => ne65_locking);
	node_ne910 : node_4 port map(clock => clock, ocupation => ocupation(4), reset => reset, R38_command => cmd_R38_ne910, R55_command => cmd_R55_ne910, R57_command => cmd_R57_ne910, R58_command => cmd_R58_ne910, R77_command => cmd_R77_ne910, state => state_ne910, locking => ne910_locking);
	node_ne912 : node_5 port map(clock => clock, ocupation => ocupation(5), reset => reset, R8_command => cmd_R8_ne912, R26_command => cmd_R26_ne912, R28_command => cmd_R28_ne912, R37_command => cmd_R37_ne912, R75_command => cmd_R75_ne912, R76_command => cmd_R76_ne912, state => state_ne912, locking => ne912_locking);
	node_ne114 : node_6 port map(clock => clock, ocupation => ocupation(6), reset => reset, R10_command => cmd_R10_ne114, R17_command => cmd_R17_ne114, R27_command => cmd_R27_ne114, R29_command => cmd_R29_ne114, R68_command => cmd_R68_ne114, R69_command => cmd_R69_ne114, R70_command => cmd_R70_ne114, R71_command => cmd_R71_ne114, R73_command => cmd_R73_ne114, state => state_ne114, locking => ne114_locking);
	node_ne288 : node_7 port map(clock => clock, ocupation => ocupation(7), reset => reset, R39_command => cmd_R39_ne288, R41_command => cmd_R41_ne288, R43_command => cmd_R43_ne288, R44_command => cmd_R44_ne288, R60_command => cmd_R60_ne288, state => state_ne288, locking => ne288_locking);
	node_ne290 : node_8 port map(clock => clock, ocupation => ocupation(8), reset => reset, R2_command => cmd_R2_ne290, R20_command => cmd_R20_ne290, R22_command => cmd_R22_ne290, R40_command => cmd_R40_ne290, R61_command => cmd_R61_ne290, R62_command => cmd_R62_ne290, state => state_ne290, locking => ne290_locking);
	node_ne292 : node_9 port map(clock => clock, ocupation => ocupation(9), reset => reset, R21_command => cmd_R21_ne292, R22_command => cmd_R22_ne292, R61_command => cmd_R61_ne292, R88_command => cmd_R88_ne292, state => state_ne292, locking => ne292_locking);
	node_ne295 : node_10 port map(clock => clock, ocupation => ocupation(10), reset => reset, R41_command => cmd_R41_ne295, R43_command => cmd_R43_ne295, R45_command => cmd_R45_ne295, R46_command => cmd_R46_ne295, state => state_ne295, locking => ne295_locking);
	node_ne297 : node_11 port map(clock => clock, ocupation => ocupation(11), reset => reset, R11_command => cmd_R11_ne297, R42_command => cmd_R42_ne297, R45_command => cmd_R45_ne297, R46_command => cmd_R46_ne297, R47_command => cmd_R47_ne297, R85_command => cmd_R85_ne297, R86_command => cmd_R86_ne297, R87_command => cmd_R87_ne297, R89_command => cmd_R89_ne297, state => state_ne297, locking => ne297_locking);
	node_ne377 : node_12 port map(clock => clock, ocupation => ocupation(12), reset => reset, R2_command => cmd_R2_ne377, R3_command => cmd_R3_ne377, R12_command => cmd_R12_ne377, R62_command => cmd_R62_ne377, state => state_ne377, locking => ne377_locking);
	node_ne384 : node_13 port map(clock => clock, ocupation => ocupation(13), reset => reset, R11_command => cmd_R11_ne384, R42_command => cmd_R42_ne384, R47_command => cmd_R47_ne384, R59_command => cmd_R59_ne384, R60_command => cmd_R60_ne384, state => state_ne384, locking => ne384_locking);
	node_ne400 : node_14 port map(clock => clock, ocupation => ocupation(14), reset => reset, R13_command => cmd_R13_ne400, R48_command => cmd_R48_ne400, R49_command => cmd_R49_ne400, R50_command => cmd_R50_ne400, R52_command => cmd_R52_ne400, R81_command => cmd_R81_ne400, R82_command => cmd_R82_ne400, R83_command => cmd_R83_ne400, R84_command => cmd_R84_ne400, state => state_ne400, locking => ne400_locking);
	node_ne404 : node_15 port map(clock => clock, ocupation => ocupation(15), reset => reset, R48_command => cmd_R48_ne404, R49_command => cmd_R49_ne404, R51_command => cmd_R51_ne404, R53_command => cmd_R53_ne404, state => state_ne404, locking => ne404_locking);
	node_ne407 : node_16 port map(clock => clock, ocupation => ocupation(16), reset => reset, R13_command => cmd_R13_ne407, R50_command => cmd_R50_ne407, R52_command => cmd_R52_ne407, R63_command => cmd_R63_ne407, R64_command => cmd_R64_ne407, state => state_ne407, locking => ne407_locking);
	node_ne421 : node_17 port map(clock => clock, ocupation => ocupation(17), reset => reset, R4_command => cmd_R4_ne421, R5_command => cmd_R5_ne421, R14_command => cmd_R14_ne421, R67_command => cmd_R67_ne421, state => state_ne421, locking => ne421_locking);
	node_ne450 : node_18 port map(clock => clock, ocupation => ocupation(18), reset => reset, R6_command => cmd_R6_ne450, R7_command => cmd_R7_ne450, R72_command => cmd_R72_ne450, R74_command => cmd_R74_ne450, state => state_ne450, locking => ne450_locking);
	node_ne465 : node_19 port map(clock => clock, ocupation => ocupation(19), reset => reset, R8_command => cmd_R8_ne465, R9_command => cmd_R9_ne465, R15_command => cmd_R15_ne465, R75_command => cmd_R75_ne465, state => state_ne465, locking => ne465_locking);
	node_ne98 : node_20 port map(clock => clock, ocupation => ocupation(20), reset => reset, R18_command => cmd_R18_ne98, R23_command => cmd_R23_ne98, R30_command => cmd_R30_ne98, R31_command => cmd_R31_ne98, R34_command => cmd_R34_ne98, R51_command => cmd_R51_ne98, R64_command => cmd_R64_ne98, state => state_ne98, locking => ne98_locking);
	node_ne99 : node_21 port map(clock => clock, ocupation => ocupation(21), reset => reset, R30_command => cmd_R30_ne99, R34_command => cmd_R34_ne99, R35_command => cmd_R35_ne99, R36_command => cmd_R36_ne99, R51_command => cmd_R51_ne99, R64_command => cmd_R64_ne99, state => state_ne99, locking => ne99_locking);
	node_ne100 : node_22 port map(clock => clock, ocupation => ocupation(22), reset => reset, R19_command => cmd_R19_ne100, R24_command => cmd_R24_ne100, R25_command => cmd_R25_ne100, R32_command => cmd_R32_ne100, R33_command => cmd_R33_ne100, state => state_ne100, locking => ne100_locking);
	node_ne101 : node_23 port map(clock => clock, ocupation => ocupation(23), reset => reset, R25_command => cmd_R25_ne101, R26_command => cmd_R26_ne101, R32_command => cmd_R32_ne101, R37_command => cmd_R37_ne101, R38_command => cmd_R38_ne101, R55_command => cmd_R55_ne101, R77_command => cmd_R77_ne101, state => state_ne101, locking => ne101_locking);
	node_ne102 : node_24 port map(clock => clock, ocupation => ocupation(24), reset => reset, R10_command => cmd_R10_ne102, R29_command => cmd_R29_ne102, state => state_ne102, locking => ne102_locking);
	node_ne104 : node_25 port map(clock => clock, ocupation => ocupation(25), reset => reset, R11_command => cmd_R11_ne104, R59_command => cmd_R59_ne104, state => state_ne104, locking => ne104_locking);
	node_ne110 : node_26 port map(clock => clock, ocupation => ocupation(26), reset => reset, R42_command => cmd_R42_ne110, R44_command => cmd_R44_ne110, R60_command => cmd_R60_ne110, state => state_ne110, locking => ne110_locking);
	node_ne111 : node_27 port map(clock => clock, ocupation => ocupation(27), reset => reset, R2_command => cmd_R2_ne111, R62_command => cmd_R62_ne111, state => state_ne111, locking => ne111_locking);
	node_ne113 : node_28 port map(clock => clock, ocupation => ocupation(28), reset => reset, R3_command => cmd_R3_ne113, R12_command => cmd_R12_ne113, state => state_ne113, locking => ne113_locking);
	node_ne122 : node_29 port map(clock => clock, ocupation => ocupation(29), reset => reset, R13_command => cmd_R13_ne122, R63_command => cmd_R63_ne122, state => state_ne122, locking => ne122_locking);
	node_ne123 : node_30 port map(clock => clock, ocupation => ocupation(30), reset => reset, R52_command => cmd_R52_ne123, R54_command => cmd_R54_ne123, R64_command => cmd_R64_ne123, state => state_ne123, locking => ne123_locking);
	node_ne124 : node_31 port map(clock => clock, ocupation => ocupation(31), reset => reset, R4_command => cmd_R4_ne124, R67_command => cmd_R67_ne124, state => state_ne124, locking => ne124_locking);
	node_ne126 : node_32 port map(clock => clock, ocupation => ocupation(32), reset => reset, R5_command => cmd_R5_ne126, R14_command => cmd_R14_ne126, state => state_ne126, locking => ne126_locking);
	node_ne127 : node_33 port map(clock => clock, ocupation => ocupation(33), reset => reset, R6_command => cmd_R6_ne127, R16_command => cmd_R16_ne127, R56_command => cmd_R56_ne127, R69_command => cmd_R69_ne127, R71_command => cmd_R71_ne127, R72_command => cmd_R72_ne127, R77_command => cmd_R77_ne127, R78_command => cmd_R78_ne127, state => state_ne127, locking => ne127_locking);
	node_ne129 : node_34 port map(clock => clock, ocupation => ocupation(34), reset => reset, R69_command => cmd_R69_ne129, R70_command => cmd_R70_ne129, R71_command => cmd_R71_ne129, R73_command => cmd_R73_ne129, state => state_ne129, locking => ne129_locking);
	node_ne130 : node_35 port map(clock => clock, ocupation => ocupation(35), reset => reset, R7_command => cmd_R7_ne130, R55_command => cmd_R55_ne130, R57_command => cmd_R57_ne130, R70_command => cmd_R70_ne130, R73_command => cmd_R73_ne130, R74_command => cmd_R74_ne130, state => state_ne130, locking => ne130_locking);
	node_ne131 : node_36 port map(clock => clock, ocupation => ocupation(36), reset => reset, R8_command => cmd_R8_ne131, R75_command => cmd_R75_ne131, state => state_ne131, locking => ne131_locking);
	node_ne132 : node_37 port map(clock => clock, ocupation => ocupation(37), reset => reset, R27_command => cmd_R27_ne132, R28_command => cmd_R28_ne132, R68_command => cmd_R68_ne132, R76_command => cmd_R76_ne132, state => state_ne132, locking => ne132_locking);
	node_ne133 : node_38 port map(clock => clock, ocupation => ocupation(38), reset => reset, R9_command => cmd_R9_ne133, R15_command => cmd_R15_ne133, state => state_ne133, locking => ne133_locking);
	node_ne134 : node_39 port map(clock => clock, ocupation => ocupation(39), reset => reset, R16_command => cmd_R16_ne134, R78_command => cmd_R78_ne134, state => state_ne134, locking => ne134_locking);
	node_ne135 : node_40 port map(clock => clock, ocupation => ocupation(40), reset => reset, R56_command => cmd_R56_ne135, R58_command => cmd_R58_ne135, R77_command => cmd_R77_ne135, state => state_ne135, locking => ne135_locking);
	node_ne992 : node_41 port map(clock => clock, ocupation => ocupation(41), reset => reset, R24_command => cmd_R24_ne992, R33_command => cmd_R33_ne992, R79_command => cmd_R79_ne992, R80_command => cmd_R80_ne992, R81_command => cmd_R81_ne992, R84_command => cmd_R84_ne992, state => state_ne992, locking => ne992_locking);
	node_ne993 : node_42 port map(clock => clock, ocupation => ocupation(42), reset => reset, R82_command => cmd_R82_ne993, R83_command => cmd_R83_ne993, state => state_ne993, locking => ne993_locking);
	node_ne994 : node_43 port map(clock => clock, ocupation => ocupation(43), reset => reset, R81_command => cmd_R81_ne994, R84_command => cmd_R84_ne994, state => state_ne994, locking => ne994_locking);
	node_ne995 : node_44 port map(clock => clock, ocupation => ocupation(44), reset => reset, R85_command => cmd_R85_ne995, R86_command => cmd_R86_ne995, state => state_ne995, locking => ne995_locking);
	node_ne996 : node_45 port map(clock => clock, ocupation => ocupation(45), reset => reset, R21_command => cmd_R21_ne996, R23_command => cmd_R23_ne996, R31_command => cmd_R31_ne996, R87_command => cmd_R87_ne996, R88_command => cmd_R88_ne996, R89_command => cmd_R89_ne996, state => state_ne996, locking => ne996_locking);
	node_ne997 : node_46 port map(clock => clock, ocupation => ocupation(46), reset => reset, R87_command => cmd_R87_ne997, R89_command => cmd_R89_ne997, state => state_ne997, locking => ne997_locking);
	route_R1 : route_0 port map(clock => clock, routeRequest => routes_i(0), reset => reset, ne991_command => cmd_R1_ne991, ne991_state => state_ne991, ne991_lock => ne991_locking, T02_state => state_T02, T02_lock => T02_locking, T02_command => cmd_R1_T02, S64_state => state_S64, routeState => routes_o(0));
	route_R2 : route_1 port map(clock => clock, routeRequest => routes_i(1), reset => reset, ne290_command => cmd_R2_ne290, ne290_state => state_ne290, ne290_lock => ne290_locking, ne377_command => cmd_R2_ne377, ne377_state => state_ne377, ne377_lock => ne377_locking, ne111_command => cmd_R2_ne111, ne111_state => state_ne111, ne111_lock => ne111_locking, D14_command => cmd_R2_D14, D14_state => state_D14, D14_lock => D14_locking, D15_command => cmd_R2_D15, D15_state => state_D15, D15_lock => D15_locking, T04_state => state_T04, T04_lock => T04_locking, T04_command => cmd_R2_T04, J35_state => state_J35, routeState => routes_o(1));
	route_R3 : route_2 port map(clock => clock, routeRequest => routes_i(2), reset => reset, ne377_command => cmd_R3_ne377, ne377_state => state_ne377, ne377_lock => ne377_locking, ne113_command => cmd_R3_ne113, ne113_state => state_ne113, ne113_lock => ne113_locking, D15_command => cmd_R3_D15, D15_state => state_D15, D15_lock => D15_locking, T04_state => state_T04, T04_lock => T04_locking, T04_command => cmd_R3_T04, T15_state => state_T15, routeState => routes_o(2));
	route_R4 : route_3 port map(clock => clock, routeRequest => routes_i(3), reset => reset, ne63_command => cmd_R4_ne63, ne63_state => state_ne63, ne63_lock => ne63_locking, ne421_command => cmd_R4_ne421, ne421_state => state_ne421, ne421_lock => ne421_locking, ne124_command => cmd_R4_ne124, ne124_state => state_ne124, ne124_lock => ne124_locking, D18_command => cmd_R4_D18, D18_state => state_D18, D18_lock => D18_locking, D19_command => cmd_R4_D19, D19_state => state_D19, D19_lock => D19_locking, T06_state => state_T06, T06_lock => T06_locking, T06_command => cmd_R4_T06, C54_state => state_C54, routeState => routes_o(3));
	route_R5 : route_4 port map(clock => clock, routeRequest => routes_i(4), reset => reset, ne421_command => cmd_R5_ne421, ne421_state => state_ne421, ne421_lock => ne421_locking, ne126_command => cmd_R5_ne126, ne126_state => state_ne126, ne126_lock => ne126_locking, D19_command => cmd_R5_D19, D19_state => state_D19, D19_lock => D19_locking, T06_state => state_T06, T06_lock => T06_locking, T06_command => cmd_R5_T06, T19_state => state_T19, routeState => routes_o(4));
	route_R6 : route_5 port map(clock => clock, routeRequest => routes_i(5), reset => reset, ne450_command => cmd_R6_ne450, ne450_state => state_ne450, ne450_lock => ne450_locking, ne127_command => cmd_R6_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, D12_command => cmd_R6_D12, D12_state => state_D12, D12_lock => D12_locking, T08_state => state_T08, T08_lock => T08_locking, T08_command => cmd_R6_T08, S117_state => state_S117, routeState => routes_o(5));
	route_R7 : route_6 port map(clock => clock, routeRequest => routes_i(6), reset => reset, ne450_command => cmd_R7_ne450, ne450_state => state_ne450, ne450_lock => ne450_locking, ne130_command => cmd_R7_ne130, ne130_state => state_ne130, ne130_lock => ne130_locking, D12_command => cmd_R7_D12, D12_state => state_D12, D12_lock => D12_locking, T08_state => state_T08, T08_lock => T08_locking, T08_command => cmd_R7_T08, C79_state => state_C79, routeState => routes_o(6));
	route_R8 : route_7 port map(clock => clock, routeRequest => routes_i(7), reset => reset, ne912_command => cmd_R8_ne912, ne912_state => state_ne912, ne912_lock => ne912_locking, ne465_command => cmd_R8_ne465, ne465_state => state_ne465, ne465_lock => ne465_locking, ne131_command => cmd_R8_ne131, ne131_state => state_ne131, ne131_lock => ne131_locking, D20_command => cmd_R8_D20, D20_state => state_D20, D20_lock => D20_locking, D21_command => cmd_R8_D21, D21_state => state_D21, D21_lock => D21_locking, T10_state => state_T10, T10_lock => T10_locking, T10_command => cmd_R8_T10, J45_state => state_J45, routeState => routes_o(7));
	route_R9 : route_8 port map(clock => clock, routeRequest => routes_i(8), reset => reset, ne465_command => cmd_R9_ne465, ne465_state => state_ne465, ne465_lock => ne465_locking, ne133_command => cmd_R9_ne133, ne133_state => state_ne133, ne133_lock => ne133_locking, D21_command => cmd_R9_D21, D21_state => state_D21, D21_lock => D21_locking, T10_state => state_T10, T10_lock => T10_locking, T10_command => cmd_R9_T10, T21_state => state_T21, routeState => routes_o(8));
	route_R10 : route_9 port map(clock => clock, routeRequest => routes_i(9), reset => reset, ne114_command => cmd_R10_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne102_command => cmd_R10_ne102, ne102_state => state_ne102, ne102_lock => ne102_locking, T12_state => state_T12, T12_lock => T12_locking, T12_command => cmd_R10_T12, S101_state => state_S101, routeState => routes_o(9));
	route_R11 : route_10 port map(clock => clock, routeRequest => routes_i(10), reset => reset, ne297_command => cmd_R11_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, ne384_command => cmd_R11_ne384, ne384_state => state_ne384, ne384_lock => ne384_locking, ne104_command => cmd_R11_ne104, ne104_state => state_ne104, ne104_lock => ne104_locking, D04_command => cmd_R11_D04, D04_state => state_D04, D04_lock => D04_locking, Sw02_command => cmd_R11_Sw02, Sw02_state => state_Sw02, Sw02_lock => Sw02_locking, T14_state => state_T14, T14_lock => T14_locking, T14_command => cmd_R11_T14, S126_state => state_S126, routeState => routes_o(10));
	route_R12 : route_11 port map(clock => clock, routeRequest => routes_i(11), reset => reset, ne377_command => cmd_R12_ne377, ne377_state => state_ne377, ne377_lock => ne377_locking, ne113_command => cmd_R12_ne113, ne113_state => state_ne113, ne113_lock => ne113_locking, D15_command => cmd_R12_D15, D15_state => state_D15, D15_lock => D15_locking, T16_state => state_T16, T16_lock => T16_locking, T16_command => cmd_R12_T16, T03_state => state_T03, routeState => routes_o(11));
	route_R13 : route_12 port map(clock => clock, routeRequest => routes_i(12), reset => reset, ne400_command => cmd_R13_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne407_command => cmd_R13_ne407, ne407_state => state_ne407, ne407_lock => ne407_locking, ne122_command => cmd_R13_ne122, ne122_state => state_ne122, ne122_lock => ne122_locking, D07_command => cmd_R13_D07, D07_state => state_D07, D07_lock => D07_locking, D16_command => cmd_R13_D16, D16_state => state_D16, D16_lock => D16_locking, T18_state => state_T18, T18_lock => T18_locking, T18_command => cmd_R13_T18, S123_state => state_S123, routeState => routes_o(12));
	route_R14 : route_13 port map(clock => clock, routeRequest => routes_i(13), reset => reset, ne421_command => cmd_R14_ne421, ne421_state => state_ne421, ne421_lock => ne421_locking, ne126_command => cmd_R14_ne126, ne126_state => state_ne126, ne126_lock => ne126_locking, D19_command => cmd_R14_D19, D19_state => state_D19, D19_lock => D19_locking, T20_state => state_T20, T20_lock => T20_locking, T20_command => cmd_R14_T20, T05_state => state_T05, routeState => routes_o(13));
	route_R15 : route_14 port map(clock => clock, routeRequest => routes_i(14), reset => reset, ne465_command => cmd_R15_ne465, ne465_state => state_ne465, ne465_lock => ne465_locking, ne133_command => cmd_R15_ne133, ne133_state => state_ne133, ne133_lock => ne133_locking, D21_command => cmd_R15_D21, D21_state => state_D21, D21_lock => D21_locking, T22_state => state_T22, T22_lock => T22_locking, T22_command => cmd_R15_T22, T09_state => state_T09, routeState => routes_o(14));
	route_R16 : route_15 port map(clock => clock, routeRequest => routes_i(15), reset => reset, ne127_command => cmd_R16_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, ne134_command => cmd_R16_ne134, ne134_state => state_ne134, ne134_lock => ne134_locking, D24_command => cmd_R16_D24, D24_state => state_D24, D24_lock => D24_locking, T24_state => state_T24, T24_lock => T24_locking, T24_command => cmd_R16_T24, S104_state => state_S104, routeState => routes_o(15));
	route_R17 : route_16 port map(clock => clock, routeRequest => routes_i(16), reset => reset, ne114_command => cmd_R17_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, L29_state => state_L29, L29_lock => L29_locking, L29_command => cmd_R17_L29, J48_state => state_J48, routeState => routes_o(16));
	route_R18 : route_17 port map(clock => clock, routeRequest => routes_i(17), reset => reset, ne98_command => cmd_R18_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, L30_state => state_L30, L30_lock => L30_locking, L30_command => cmd_R18_L30, X50_state => state_X50, routeState => routes_o(17));
	route_R19 : route_18 port map(clock => clock, routeRequest => routes_i(18), reset => reset, ne100_command => cmd_R19_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, L31_state => state_L31, L31_lock => L31_locking, L31_command => cmd_R19_L31, X52_state => state_X52, routeState => routes_o(18));
	route_R20 : route_19 port map(clock => clock, routeRequest => routes_i(19), reset => reset, ne991_command => cmd_R20_ne991, ne991_state => state_ne991, ne991_lock => ne991_locking, ne290_command => cmd_R20_ne290, ne290_state => state_ne290, ne290_lock => ne290_locking, D01_command => cmd_R20_D01, D01_state => state_D01, D01_lock => D01_locking, J35_state => state_J35, J35_lock => J35_locking, J35_command => cmd_R20_J35, T01_state => state_T01, routeState => routes_o(19));
	route_R21 : route_20 port map(clock => clock, routeRequest => routes_i(20), reset => reset, ne292_command => cmd_R21_ne292, ne292_state => state_ne292, ne292_lock => ne292_locking, ne996_command => cmd_R21_ne996, ne996_state => state_ne996, ne996_lock => ne996_locking, Sw04_command => cmd_R21_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, J36_state => state_J36, J36_lock => J36_locking, J36_command => cmd_R21_J36, J38_state => state_J38, routeState => routes_o(20));
	route_R22 : route_21 port map(clock => clock, routeRequest => routes_i(21), reset => reset, ne290_command => cmd_R22_ne290, ne290_state => state_ne290, ne290_lock => ne290_locking, ne292_command => cmd_R22_ne292, ne292_state => state_ne292, ne292_lock => ne292_locking, D14_command => cmd_R22_D14, D14_state => state_D14, D14_lock => D14_locking, J37_state => state_J37, J37_lock => J37_locking, J37_command => cmd_R22_J37, J35_state => state_J35, routeState => routes_o(21));
	route_R23 : route_22 port map(clock => clock, routeRequest => routes_i(22), reset => reset, ne98_command => cmd_R23_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne996_command => cmd_R23_ne996, ne996_state => state_ne996, ne996_lock => ne996_locking, J38_state => state_J38, J38_lock => J38_locking, J38_command => cmd_R23_J38, L30_state => state_L30, routeState => routes_o(22));
	route_R24 : route_23 port map(clock => clock, routeRequest => routes_i(23), reset => reset, ne100_command => cmd_R24_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne992_command => cmd_R24_ne992, ne992_state => state_ne992, ne992_lock => ne992_locking, J40_state => state_J40, J40_lock => J40_locking, J40_command => cmd_R24_J40, L31_state => state_L31, routeState => routes_o(23));
	route_R25 : route_24 port map(clock => clock, routeRequest => routes_i(24), reset => reset, ne100_command => cmd_R25_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne101_command => cmd_R25_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, J43_state => state_J43, J43_lock => J43_locking, J43_command => cmd_R25_J43, X53_state => state_X53, routeState => routes_o(24));
	route_R26 : route_25 port map(clock => clock, routeRequest => routes_i(25), reset => reset, ne912_command => cmd_R26_ne912, ne912_state => state_ne912, ne912_lock => ne912_locking, ne101_command => cmd_R26_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, D09_command => cmd_R26_D09, D09_state => state_D09, D09_lock => D09_locking, J45_state => state_J45, J45_lock => J45_locking, J45_command => cmd_R26_J45, J43_state => state_J43, routeState => routes_o(25));
	route_R27 : route_26 port map(clock => clock, routeRequest => routes_i(26), reset => reset, ne114_command => cmd_R27_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne132_command => cmd_R27_ne132, ne132_state => state_ne132, ne132_lock => ne132_locking, D23_command => cmd_R27_D23, D23_state => state_D23, D23_lock => D23_locking, J46_state => state_J46, J46_lock => J46_locking, J46_command => cmd_R27_J46, L29_state => state_L29, routeState => routes_o(26));
	route_R28 : route_27 port map(clock => clock, routeRequest => routes_i(27), reset => reset, ne912_command => cmd_R28_ne912, ne912_state => state_ne912, ne912_lock => ne912_locking, ne132_command => cmd_R28_ne132, ne132_state => state_ne132, ne132_lock => ne132_locking, D20_command => cmd_R28_D20, D20_state => state_D20, D20_lock => D20_locking, J47_state => state_J47, J47_lock => J47_locking, J47_command => cmd_R28_J47, J45_state => state_J45, routeState => routes_o(27));
	route_R29 : route_28 port map(clock => clock, routeRequest => routes_i(28), reset => reset, ne114_command => cmd_R29_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne102_command => cmd_R29_ne102, ne102_state => state_ne102, ne102_lock => ne102_locking, J48_state => state_J48, J48_lock => J48_locking, J48_command => cmd_R29_J48, T11_state => state_T11, routeState => routes_o(28));
	route_R30 : route_29 port map(clock => clock, routeRequest => routes_i(29), reset => reset, ne98_command => cmd_R30_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne99_command => cmd_R30_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, Lc01_command => cmd_R30_Lc01, Lc01_state => state_Lc01, Lc01_lock => Lc01_locking, X50_state => state_X50, X50_lock => X50_locking, X50_command => cmd_R30_X50, S55_state => state_S55, routeState => routes_o(29));
	route_R31 : route_30 port map(clock => clock, routeRequest => routes_i(30), reset => reset, ne98_command => cmd_R31_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne996_command => cmd_R31_ne996, ne996_state => state_ne996, ne996_lock => ne996_locking, Lc01_command => cmd_R31_Lc01, Lc01_state => state_Lc01, Lc01_lock => Lc01_locking, X51_state => state_X51, X51_lock => X51_locking, X51_command => cmd_R31_X51, S129_state => state_S129, routeState => routes_o(30));
	route_R32 : route_31 port map(clock => clock, routeRequest => routes_i(31), reset => reset, ne100_command => cmd_R32_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne101_command => cmd_R32_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, Lc04_command => cmd_R32_Lc04, Lc04_state => state_Lc04, Lc04_lock => Lc04_locking, X52_state => state_X52, X52_lock => X52_locking, X52_command => cmd_R32_X52, S59_state => state_S59, routeState => routes_o(31));
	route_R33 : route_32 port map(clock => clock, routeRequest => routes_i(32), reset => reset, ne100_command => cmd_R33_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne992_command => cmd_R33_ne992, ne992_state => state_ne992, ne992_lock => ne992_locking, Lc04_command => cmd_R33_Lc04, Lc04_state => state_Lc04, Lc04_lock => Lc04_locking, X53_state => state_X53, X53_lock => X53_locking, X53_command => cmd_R33_X53, S120_state => state_S120, routeState => routes_o(32));
	route_R34 : route_33 port map(clock => clock, routeRequest => routes_i(33), reset => reset, ne63_command => cmd_R34_ne63, ne63_state => state_ne63, ne63_lock => ne63_locking, ne98_command => cmd_R34_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne99_command => cmd_R34_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, D05_command => cmd_R34_D05, D05_state => state_D05, D05_lock => D05_locking, C54_state => state_C54, C54_lock => C54_locking, C54_command => cmd_R34_C54, X51_state => state_X51, routeState => routes_o(33));
	route_R35 : route_34 port map(clock => clock, routeRequest => routes_i(34), reset => reset, ne61_command => cmd_R35_ne61, ne61_state => state_ne61, ne61_lock => ne61_locking, ne99_command => cmd_R35_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, D05_command => cmd_R35_D05, D05_state => state_D05, D05_lock => D05_locking, S55_state => state_S55, S55_lock => S55_locking, S55_command => cmd_R35_S55, S78_state => state_S78, routeState => routes_o(34));
	route_R36 : route_35 port map(clock => clock, routeRequest => routes_i(35), reset => reset, ne63_command => cmd_R36_ne63, ne63_state => state_ne63, ne63_lock => ne63_locking, ne99_command => cmd_R36_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, D05_command => cmd_R36_D05, D05_state => state_D05, D05_lock => D05_locking, S55_state => state_S55, S55_lock => S55_locking, S55_command => cmd_R36_S55, S95_state => state_S95, routeState => routes_o(35));
	route_R37 : route_36 port map(clock => clock, routeRequest => routes_i(36), reset => reset, ne912_command => cmd_R37_ne912, ne912_state => state_ne912, ne912_lock => ne912_locking, ne101_command => cmd_R37_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, D09_command => cmd_R37_D09, D09_state => state_D09, D09_lock => D09_locking, S59_state => state_S59, S59_lock => S59_locking, S59_command => cmd_R37_S59, S110_state => state_S110, routeState => routes_o(36));
	route_R38 : route_37 port map(clock => clock, routeRequest => routes_i(37), reset => reset, ne910_command => cmd_R38_ne910, ne910_state => state_ne910, ne910_lock => ne910_locking, ne101_command => cmd_R38_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, D09_command => cmd_R38_D09, D09_state => state_D09, D09_lock => D09_locking, S59_state => state_S59, S59_lock => S59_locking, S59_command => cmd_R38_S59, S81_state => state_S81, routeState => routes_o(37));
	route_R39 : route_38 port map(clock => clock, routeRequest => routes_i(38), reset => reset, ne991_command => cmd_R39_ne991, ne991_state => state_ne991, ne991_lock => ne991_locking, ne288_command => cmd_R39_ne288, ne288_state => state_ne288, ne288_lock => ne288_locking, D01_command => cmd_R39_D01, D01_state => state_D01, D01_lock => D01_locking, S64_state => state_S64, S64_lock => S64_locking, S64_command => cmd_R39_S64, S69_state => state_S69, routeState => routes_o(38));
	route_R40 : route_39 port map(clock => clock, routeRequest => routes_i(39), reset => reset, ne991_command => cmd_R40_ne991, ne991_state => state_ne991, ne991_lock => ne991_locking, ne290_command => cmd_R40_ne290, ne290_state => state_ne290, ne290_lock => ne290_locking, D01_command => cmd_R40_D01, D01_state => state_D01, D01_lock => D01_locking, S64_state => state_S64, S64_lock => S64_locking, S64_command => cmd_R40_S64, S86_state => state_S86, routeState => routes_o(39));
	route_R41 : route_40 port map(clock => clock, routeRequest => routes_i(40), reset => reset, ne991_command => cmd_R41_ne991, ne991_state => state_ne991, ne991_lock => ne991_locking, ne288_command => cmd_R41_ne288, ne288_state => state_ne288, ne288_lock => ne288_locking, ne295_command => cmd_R41_ne295, ne295_state => state_ne295, ne295_lock => ne295_locking, D01_command => cmd_R41_D01, D01_state => state_D01, D01_lock => D01_locking, D03_command => cmd_R41_D03, D03_state => state_D03, D03_lock => D03_locking, C67_state => state_C67, C67_lock => C67_locking, C67_command => cmd_R41_C67, T01_state => state_T01, routeState => routes_o(40));
	route_R42 : route_41 port map(clock => clock, routeRequest => routes_i(41), reset => reset, ne297_command => cmd_R42_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, ne384_command => cmd_R42_ne384, ne384_state => state_ne384, ne384_lock => ne384_locking, ne110_command => cmd_R42_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, D04_command => cmd_R42_D04, D04_state => state_D04, D04_lock => D04_locking, Sw02_command => cmd_R42_Sw02, Sw02_state => state_Sw02, Sw02_lock => Sw02_locking, B68_state => state_B68, B68_lock => B68_locking, B68_command => cmd_R42_B68, S126_state => state_S126, routeState => routes_o(41));
	route_R43 : route_42 port map(clock => clock, routeRequest => routes_i(42), reset => reset, ne288_command => cmd_R43_ne288, ne288_state => state_ne288, ne288_lock => ne288_locking, ne295_command => cmd_R43_ne295, ne295_state => state_ne295, ne295_lock => ne295_locking, D03_command => cmd_R43_D03, D03_state => state_D03, D03_lock => D03_locking, S69_state => state_S69, S69_lock => S69_locking, S69_command => cmd_R43_S69, C70_state => state_C70, routeState => routes_o(42));
	route_R44 : route_43 port map(clock => clock, routeRequest => routes_i(43), reset => reset, ne288_command => cmd_R44_ne288, ne288_state => state_ne288, ne288_lock => ne288_locking, ne110_command => cmd_R44_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, D03_command => cmd_R44_D03, D03_state => state_D03, D03_lock => D03_locking, S69_state => state_S69, S69_lock => S69_locking, S69_command => cmd_R44_S69, B68_state => state_B68, routeState => routes_o(43));
	route_R45 : route_44 port map(clock => clock, routeRequest => routes_i(44), reset => reset, ne295_command => cmd_R45_ne295, ne295_state => state_ne295, ne295_lock => ne295_locking, ne297_command => cmd_R45_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, D04_command => cmd_R45_D04, D04_state => state_D04, D04_lock => D04_locking, C70_state => state_C70, C70_lock => C70_locking, C70_command => cmd_R45_C70, S126_state => state_S126, routeState => routes_o(44));
	route_R46 : route_45 port map(clock => clock, routeRequest => routes_i(45), reset => reset, ne295_command => cmd_R46_ne295, ne295_state => state_ne295, ne295_lock => ne295_locking, ne297_command => cmd_R46_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, D04_command => cmd_R46_D04, D04_state => state_D04, D04_lock => D04_locking, S71_state => state_S71, S71_lock => S71_locking, S71_command => cmd_R46_S71, C67_state => state_C67, routeState => routes_o(45));
	route_R47 : route_46 port map(clock => clock, routeRequest => routes_i(46), reset => reset, ne297_command => cmd_R47_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, ne384_command => cmd_R47_ne384, ne384_state => state_ne384, ne384_lock => ne384_locking, D04_command => cmd_R47_D04, D04_state => state_D04, D04_lock => D04_locking, S71_state => state_S71, S71_lock => S71_locking, S71_command => cmd_R47_S71, S84_state => state_S84, routeState => routes_o(46));
	route_R48 : route_47 port map(clock => clock, routeRequest => routes_i(47), reset => reset, ne400_command => cmd_R48_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne404_command => cmd_R48_ne404, ne404_state => state_ne404, ne404_lock => ne404_locking, D07_command => cmd_R48_D07, D07_state => state_D07, D07_lock => D07_locking, C73_state => state_C73, C73_lock => C73_locking, C73_command => cmd_R48_C73, S123_state => state_S123, routeState => routes_o(47));
	route_R49 : route_48 port map(clock => clock, routeRequest => routes_i(48), reset => reset, ne400_command => cmd_R49_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne404_command => cmd_R49_ne404, ne404_state => state_ne404, ne404_lock => ne404_locking, D07_command => cmd_R49_D07, D07_state => state_D07, D07_lock => D07_locking, S74_state => state_S74, S74_lock => S74_locking, S74_command => cmd_R49_S74, C76_state => state_C76, routeState => routes_o(48));
	route_R50 : route_49 port map(clock => clock, routeRequest => routes_i(49), reset => reset, ne400_command => cmd_R50_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne407_command => cmd_R50_ne407, ne407_state => state_ne407, ne407_lock => ne407_locking, D07_command => cmd_R50_D07, D07_state => state_D07, D07_lock => D07_locking, S74_state => state_S74, S74_lock => S74_locking, S74_command => cmd_R50_S74, S93_state => state_S93, routeState => routes_o(49));
	route_R51 : route_50 port map(clock => clock, routeRequest => routes_i(50), reset => reset, ne61_command => cmd_R51_ne61, ne61_state => state_ne61, ne61_lock => ne61_locking, ne404_command => cmd_R51_ne404, ne404_state => state_ne404, ne404_lock => ne404_locking, ne98_command => cmd_R51_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne99_command => cmd_R51_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, D05_command => cmd_R51_D05, D05_state => state_D05, D05_lock => D05_locking, D08_command => cmd_R51_D08, D08_state => state_D08, D08_lock => D08_locking, C76_state => state_C76, C76_lock => C76_locking, C76_command => cmd_R51_C76, X51_state => state_X51, routeState => routes_o(50));
	route_R52 : route_51 port map(clock => clock, routeRequest => routes_i(51), reset => reset, ne400_command => cmd_R52_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne407_command => cmd_R52_ne407, ne407_state => state_ne407, ne407_lock => ne407_locking, ne123_command => cmd_R52_ne123, ne123_state => state_ne123, ne123_lock => ne123_locking, D07_command => cmd_R52_D07, D07_state => state_D07, D07_lock => D07_locking, D16_command => cmd_R52_D16, D16_state => state_D16, D16_lock => D16_locking, B77_state => state_B77, B77_lock => B77_locking, B77_command => cmd_R52_B77, S123_state => state_S123, routeState => routes_o(51));
	route_R53 : route_52 port map(clock => clock, routeRequest => routes_i(52), reset => reset, ne61_command => cmd_R53_ne61, ne61_state => state_ne61, ne61_lock => ne61_locking, ne404_command => cmd_R53_ne404, ne404_state => state_ne404, ne404_lock => ne404_locking, D08_command => cmd_R53_D08, D08_state => state_D08, D08_lock => D08_locking, S78_state => state_S78, S78_lock => S78_locking, S78_command => cmd_R53_S78, C73_state => state_C73, routeState => routes_o(52));
	route_R54 : route_53 port map(clock => clock, routeRequest => routes_i(53), reset => reset, ne61_command => cmd_R54_ne61, ne61_state => state_ne61, ne61_lock => ne61_locking, ne123_command => cmd_R54_ne123, ne123_state => state_ne123, ne123_lock => ne123_locking, D08_command => cmd_R54_D08, D08_state => state_D08, D08_lock => D08_locking, S78_state => state_S78, S78_lock => S78_locking, S78_command => cmd_R54_S78, B77_state => state_B77, routeState => routes_o(53));
	route_R55 : route_54 port map(clock => clock, routeRequest => routes_i(54), reset => reset, ne910_command => cmd_R55_ne910, ne910_state => state_ne910, ne910_lock => ne910_locking, ne101_command => cmd_R55_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, ne130_command => cmd_R55_ne130, ne130_state => state_ne130, ne130_lock => ne130_locking, D09_command => cmd_R55_D09, D09_state => state_D09, D09_lock => D09_locking, D10_command => cmd_R55_D10, D10_state => state_D10, D10_lock => D10_locking, C79_state => state_C79, C79_lock => C79_locking, C79_command => cmd_R55_C79, J43_state => state_J43, routeState => routes_o(54));
	route_R56 : route_55 port map(clock => clock, routeRequest => routes_i(55), reset => reset, ne127_command => cmd_R56_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, ne135_command => cmd_R56_ne135, ne135_state => state_ne135, ne135_lock => ne135_locking, D24_command => cmd_R56_D24, D24_state => state_D24, D24_lock => D24_locking, B80_state => state_B80, B80_lock => B80_locking, B80_command => cmd_R56_B80, S104_state => state_S104, routeState => routes_o(55));
	route_R57 : route_56 port map(clock => clock, routeRequest => routes_i(56), reset => reset, ne910_command => cmd_R57_ne910, ne910_state => state_ne910, ne910_lock => ne910_locking, ne130_command => cmd_R57_ne130, ne130_state => state_ne130, ne130_lock => ne130_locking, D10_command => cmd_R57_D10, D10_state => state_D10, D10_lock => D10_locking, S81_state => state_S81, S81_lock => S81_locking, S81_command => cmd_R57_S81, S107_state => state_S107, routeState => routes_o(56));
	route_R58 : route_57 port map(clock => clock, routeRequest => routes_i(57), reset => reset, ne910_command => cmd_R58_ne910, ne910_state => state_ne910, ne910_lock => ne910_locking, ne135_command => cmd_R58_ne135, ne135_state => state_ne135, ne135_lock => ne135_locking, D10_command => cmd_R58_D10, D10_state => state_D10, D10_lock => D10_locking, S81_state => state_S81, S81_lock => S81_locking, S81_command => cmd_R58_S81, B80_state => state_B80, routeState => routes_o(57));
	route_R59 : route_58 port map(clock => clock, routeRequest => routes_i(58), reset => reset, ne384_command => cmd_R59_ne384, ne384_state => state_ne384, ne384_lock => ne384_locking, ne104_command => cmd_R59_ne104, ne104_state => state_ne104, ne104_lock => ne104_locking, Sw02_command => cmd_R59_Sw02, Sw02_state => state_Sw02, Sw02_lock => Sw02_locking, S84_state => state_S84, S84_lock => S84_locking, S84_command => cmd_R59_S84, T13_state => state_T13, routeState => routes_o(58));
	route_R60 : route_59 port map(clock => clock, routeRequest => routes_i(59), reset => reset, ne991_command => cmd_R60_ne991, ne991_state => state_ne991, ne991_lock => ne991_locking, ne288_command => cmd_R60_ne288, ne288_state => state_ne288, ne288_lock => ne288_locking, ne384_command => cmd_R60_ne384, ne384_state => state_ne384, ne384_lock => ne384_locking, ne110_command => cmd_R60_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, D01_command => cmd_R60_D01, D01_state => state_D01, D01_lock => D01_locking, D03_command => cmd_R60_D03, D03_state => state_D03, D03_lock => D03_locking, Sw02_command => cmd_R60_Sw02, Sw02_state => state_Sw02, Sw02_lock => Sw02_locking, S84_state => state_S84, S84_lock => S84_locking, S84_command => cmd_R60_S84, T01_state => state_T01, routeState => routes_o(59));
	route_R61 : route_60 port map(clock => clock, routeRequest => routes_i(60), reset => reset, ne290_command => cmd_R61_ne290, ne290_state => state_ne290, ne290_lock => ne290_locking, ne292_command => cmd_R61_ne292, ne292_state => state_ne292, ne292_lock => ne292_locking, D14_command => cmd_R61_D14, D14_state => state_D14, D14_lock => D14_locking, S86_state => state_S86, S86_lock => S86_locking, S86_command => cmd_R61_S86, J36_state => state_J36, routeState => routes_o(60));
	route_R62 : route_61 port map(clock => clock, routeRequest => routes_i(61), reset => reset, ne290_command => cmd_R62_ne290, ne290_state => state_ne290, ne290_lock => ne290_locking, ne377_command => cmd_R62_ne377, ne377_state => state_ne377, ne377_lock => ne377_locking, ne111_command => cmd_R62_ne111, ne111_state => state_ne111, ne111_lock => ne111_locking, D14_command => cmd_R62_D14, D14_state => state_D14, D14_lock => D14_locking, D15_command => cmd_R62_D15, D15_state => state_D15, D15_lock => D15_locking, S86_state => state_S86, S86_lock => S86_locking, S86_command => cmd_R62_S86, T03_state => state_T03, routeState => routes_o(61));
	route_R63 : route_62 port map(clock => clock, routeRequest => routes_i(62), reset => reset, ne407_command => cmd_R63_ne407, ne407_state => state_ne407, ne407_lock => ne407_locking, ne122_command => cmd_R63_ne122, ne122_state => state_ne122, ne122_lock => ne122_locking, D16_command => cmd_R63_D16, D16_state => state_D16, D16_lock => D16_locking, S93_state => state_S93, S93_lock => S93_locking, S93_command => cmd_R63_S93, T17_state => state_T17, routeState => routes_o(62));
	route_R64 : route_63 port map(clock => clock, routeRequest => routes_i(63), reset => reset, ne61_command => cmd_R64_ne61, ne61_state => state_ne61, ne61_lock => ne61_locking, ne407_command => cmd_R64_ne407, ne407_state => state_ne407, ne407_lock => ne407_locking, ne98_command => cmd_R64_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne99_command => cmd_R64_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, ne123_command => cmd_R64_ne123, ne123_state => state_ne123, ne123_lock => ne123_locking, D05_command => cmd_R64_D05, D05_state => state_D05, D05_lock => D05_locking, D08_command => cmd_R64_D08, D08_state => state_D08, D08_lock => D08_locking, D16_command => cmd_R64_D16, D16_state => state_D16, D16_lock => D16_locking, S93_state => state_S93, S93_lock => S93_locking, S93_command => cmd_R64_S93, X51_state => state_X51, routeState => routes_o(63));
	route_R65 : route_64 port map(clock => clock, routeRequest => routes_i(64), reset => reset, ne63_command => cmd_R65_ne63, ne63_state => state_ne63, ne63_lock => ne63_locking, ne65_command => cmd_R65_ne65, ne65_state => state_ne65, ne65_lock => ne65_locking, D18_command => cmd_R65_D18, D18_state => state_D18, D18_lock => D18_locking, C94_state => state_C94, C94_lock => C94_locking, C94_command => cmd_R65_C94, C54_state => state_C54, routeState => routes_o(64));
	route_R66 : route_65 port map(clock => clock, routeRequest => routes_i(65), reset => reset, ne63_command => cmd_R66_ne63, ne63_state => state_ne63, ne63_lock => ne63_locking, ne65_command => cmd_R66_ne65, ne65_state => state_ne65, ne65_lock => ne65_locking, D18_command => cmd_R66_D18, D18_state => state_D18, D18_lock => D18_locking, S95_state => state_S95, S95_lock => S95_locking, S95_command => cmd_R66_S95, C119_state => state_C119, routeState => routes_o(65));
	route_R67 : route_66 port map(clock => clock, routeRequest => routes_i(66), reset => reset, ne63_command => cmd_R67_ne63, ne63_state => state_ne63, ne63_lock => ne63_locking, ne421_command => cmd_R67_ne421, ne421_state => state_ne421, ne421_lock => ne421_locking, ne124_command => cmd_R67_ne124, ne124_state => state_ne124, ne124_lock => ne124_locking, D18_command => cmd_R67_D18, D18_state => state_D18, D18_lock => D18_locking, D19_command => cmd_R67_D19, D19_state => state_D19, D19_lock => D19_locking, S95_state => state_S95, S95_lock => S95_locking, S95_command => cmd_R67_S95, T05_state => state_T05, routeState => routes_o(66));
	route_R68 : route_67 port map(clock => clock, routeRequest => routes_i(67), reset => reset, ne114_command => cmd_R68_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne132_command => cmd_R68_ne132, ne132_state => state_ne132, ne132_lock => ne132_locking, D23_command => cmd_R68_D23, D23_state => state_D23, D23_lock => D23_locking, S101_state => state_S101, S101_lock => S101_locking, S101_command => cmd_R68_S101, J47_state => state_J47, routeState => routes_o(67));
	route_R69 : route_68 port map(clock => clock, routeRequest => routes_i(68), reset => reset, ne114_command => cmd_R69_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne127_command => cmd_R69_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, ne129_command => cmd_R69_ne129, ne129_state => state_ne129, ne129_lock => ne129_locking, D23_command => cmd_R69_D23, D23_state => state_D23, D23_lock => D23_locking, D12_command => cmd_R69_D12, D12_state => state_D12, D12_lock => D12_locking, S101_state => state_S101, S101_lock => S101_locking, S101_command => cmd_R69_S101, S117_state => state_S117, routeState => routes_o(68));
	route_R70 : route_69 port map(clock => clock, routeRequest => routes_i(69), reset => reset, ne114_command => cmd_R70_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne129_command => cmd_R70_ne129, ne129_state => state_ne129, ne129_lock => ne129_locking, ne130_command => cmd_R70_ne130, ne130_state => state_ne130, ne130_lock => ne130_locking, D23_command => cmd_R70_D23, D23_state => state_D23, D23_lock => D23_locking, D12_command => cmd_R70_D12, D12_state => state_D12, D12_lock => D12_locking, S101_state => state_S101, S101_lock => S101_locking, S101_command => cmd_R70_S101, C79_state => state_C79, routeState => routes_o(69));
	route_R71 : route_70 port map(clock => clock, routeRequest => routes_i(70), reset => reset, ne114_command => cmd_R71_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne127_command => cmd_R71_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, ne129_command => cmd_R71_ne129, ne129_state => state_ne129, ne129_lock => ne129_locking, D23_command => cmd_R71_D23, D23_state => state_D23, D23_lock => D23_locking, D12_command => cmd_R71_D12, D12_state => state_D12, D12_lock => D12_locking, S104_state => state_S104, S104_lock => S104_locking, S104_command => cmd_R71_S104, L29_state => state_L29, routeState => routes_o(70));
	route_R72 : route_71 port map(clock => clock, routeRequest => routes_i(71), reset => reset, ne450_command => cmd_R72_ne450, ne450_state => state_ne450, ne450_lock => ne450_locking, ne127_command => cmd_R72_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, D12_command => cmd_R72_D12, D12_state => state_D12, D12_lock => D12_locking, S104_state => state_S104, S104_lock => S104_locking, S104_command => cmd_R72_S104, T07_state => state_T07, routeState => routes_o(71));
	route_R73 : route_72 port map(clock => clock, routeRequest => routes_i(72), reset => reset, ne114_command => cmd_R73_ne114, ne114_state => state_ne114, ne114_lock => ne114_locking, ne129_command => cmd_R73_ne129, ne129_state => state_ne129, ne129_lock => ne129_locking, ne130_command => cmd_R73_ne130, ne130_state => state_ne130, ne130_lock => ne130_locking, D23_command => cmd_R73_D23, D23_state => state_D23, D23_lock => D23_locking, D12_command => cmd_R73_D12, D12_state => state_D12, D12_lock => D12_locking, S107_state => state_S107, S107_lock => S107_locking, S107_command => cmd_R73_S107, L29_state => state_L29, routeState => routes_o(72));
	route_R74 : route_73 port map(clock => clock, routeRequest => routes_i(73), reset => reset, ne450_command => cmd_R74_ne450, ne450_state => state_ne450, ne450_lock => ne450_locking, ne130_command => cmd_R74_ne130, ne130_state => state_ne130, ne130_lock => ne130_locking, D12_command => cmd_R74_D12, D12_state => state_D12, D12_lock => D12_locking, S107_state => state_S107, S107_lock => S107_locking, S107_command => cmd_R74_S107, T07_state => state_T07, routeState => routes_o(73));
	route_R75 : route_74 port map(clock => clock, routeRequest => routes_i(74), reset => reset, ne912_command => cmd_R75_ne912, ne912_state => state_ne912, ne912_lock => ne912_locking, ne465_command => cmd_R75_ne465, ne465_state => state_ne465, ne465_lock => ne465_locking, ne131_command => cmd_R75_ne131, ne131_state => state_ne131, ne131_lock => ne131_locking, D20_command => cmd_R75_D20, D20_state => state_D20, D20_lock => D20_locking, D21_command => cmd_R75_D21, D21_state => state_D21, D21_lock => D21_locking, S110_state => state_S110, S110_lock => S110_locking, S110_command => cmd_R75_S110, T09_state => state_T09, routeState => routes_o(74));
	route_R76 : route_75 port map(clock => clock, routeRequest => routes_i(75), reset => reset, ne912_command => cmd_R76_ne912, ne912_state => state_ne912, ne912_lock => ne912_locking, ne132_command => cmd_R76_ne132, ne132_state => state_ne132, ne132_lock => ne132_locking, D20_command => cmd_R76_D20, D20_state => state_D20, D20_lock => D20_locking, S110_state => state_S110, S110_lock => S110_locking, S110_command => cmd_R76_S110, J46_state => state_J46, routeState => routes_o(75));
	route_R77 : route_76 port map(clock => clock, routeRequest => routes_i(76), reset => reset, ne910_command => cmd_R77_ne910, ne910_state => state_ne910, ne910_lock => ne910_locking, ne101_command => cmd_R77_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, ne127_command => cmd_R77_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, ne135_command => cmd_R77_ne135, ne135_state => state_ne135, ne135_lock => ne135_locking, D09_command => cmd_R77_D09, D09_state => state_D09, D09_lock => D09_locking, D10_command => cmd_R77_D10, D10_state => state_D10, D10_lock => D10_locking, D24_command => cmd_R77_D24, D24_state => state_D24, D24_lock => D24_locking, S117_state => state_S117, S117_lock => S117_locking, S117_command => cmd_R77_S117, J43_state => state_J43, routeState => routes_o(76));
	route_R78 : route_77 port map(clock => clock, routeRequest => routes_i(77), reset => reset, ne127_command => cmd_R78_ne127, ne127_state => state_ne127, ne127_lock => ne127_locking, ne134_command => cmd_R78_ne134, ne134_state => state_ne134, ne134_lock => ne134_locking, D24_command => cmd_R78_D24, D24_state => state_D24, D24_lock => D24_locking, S117_state => state_S117, S117_lock => S117_locking, S117_command => cmd_R78_S117, T23_state => state_T23, routeState => routes_o(77));
	route_R79 : route_78 port map(clock => clock, routeRequest => routes_i(78), reset => reset, ne65_command => cmd_R79_ne65, ne65_state => state_ne65, ne65_lock => ne65_locking, ne992_command => cmd_R79_ne992, ne992_state => state_ne992, ne992_lock => ne992_locking, Sw01_command => cmd_R79_Sw01, Sw01_state => state_Sw01, Sw01_lock => Sw01_locking, C119_state => state_C119, C119_lock => C119_locking, C119_command => cmd_R79_C119, J40_state => state_J40, routeState => routes_o(78));
	route_R80 : route_79 port map(clock => clock, routeRequest => routes_i(79), reset => reset, ne65_command => cmd_R80_ne65, ne65_state => state_ne65, ne65_lock => ne65_locking, ne992_command => cmd_R80_ne992, ne992_state => state_ne992, ne992_lock => ne992_locking, Sw01_command => cmd_R80_Sw01, Sw01_state => state_Sw01, Sw01_lock => Sw01_locking, S120_state => state_S120, S120_lock => S120_locking, S120_command => cmd_R80_S120, C94_state => state_C94, routeState => routes_o(79));
	route_R81 : route_80 port map(clock => clock, routeRequest => routes_i(80), reset => reset, ne400_command => cmd_R81_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne992_command => cmd_R81_ne992, ne992_state => state_ne992, ne992_lock => ne992_locking, ne994_command => cmd_R81_ne994, ne994_state => state_ne994, ne994_lock => ne994_locking, Sw01_command => cmd_R81_Sw01, Sw01_state => state_Sw01, Sw01_lock => Sw01_locking, Sw05_command => cmd_R81_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, S120_state => state_S120, S120_lock => S120_locking, S120_command => cmd_R81_S120, S74_state => state_S74, routeState => routes_o(80));
	route_R82 : route_81 port map(clock => clock, routeRequest => routes_i(81), reset => reset, ne400_command => cmd_R82_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne993_command => cmd_R82_ne993, ne993_state => state_ne993, ne993_lock => ne993_locking, Sw05_command => cmd_R82_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, C122_state => state_C122, C122_lock => C122_locking, C122_command => cmd_R82_C122, S74_state => state_S74, routeState => routes_o(81));
	route_R83 : route_82 port map(clock => clock, routeRequest => routes_i(82), reset => reset, ne400_command => cmd_R83_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne993_command => cmd_R83_ne993, ne993_state => state_ne993, ne993_lock => ne993_locking, Sw05_command => cmd_R83_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, S123_state => state_S123, S123_lock => S123_locking, S123_command => cmd_R83_S123, T25_state => state_T25, routeState => routes_o(82));
	route_R84 : route_83 port map(clock => clock, routeRequest => routes_i(83), reset => reset, ne400_command => cmd_R84_ne400, ne400_state => state_ne400, ne400_lock => ne400_locking, ne992_command => cmd_R84_ne992, ne992_state => state_ne992, ne992_lock => ne992_locking, ne994_command => cmd_R84_ne994, ne994_state => state_ne994, ne994_lock => ne994_locking, Sw01_command => cmd_R84_Sw01, Sw01_state => state_Sw01, Sw01_lock => Sw01_locking, Sw05_command => cmd_R84_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, S123_state => state_S123, S123_lock => S123_locking, S123_command => cmd_R84_S123, J40_state => state_J40, routeState => routes_o(83));
	route_R85 : route_84 port map(clock => clock, routeRequest => routes_i(84), reset => reset, ne297_command => cmd_R85_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, ne995_command => cmd_R85_ne995, ne995_state => state_ne995, ne995_lock => ne995_locking, Sw03_command => cmd_R85_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, C125_state => state_C125, C125_lock => C125_locking, C125_command => cmd_R85_C125, S71_state => state_S71, routeState => routes_o(84));
	route_R86 : route_85 port map(clock => clock, routeRequest => routes_i(85), reset => reset, ne297_command => cmd_R86_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, ne995_command => cmd_R86_ne995, ne995_state => state_ne995, ne995_lock => ne995_locking, Sw03_command => cmd_R86_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, S126_state => state_S126, S126_lock => S126_locking, S126_command => cmd_R86_S126, T27_state => state_T27, routeState => routes_o(85));
	route_R87 : route_86 port map(clock => clock, routeRequest => routes_i(86), reset => reset, ne297_command => cmd_R87_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, ne996_command => cmd_R87_ne996, ne996_state => state_ne996, ne996_lock => ne996_locking, ne997_command => cmd_R87_ne997, ne997_state => state_ne997, ne997_lock => ne997_locking, Sw03_command => cmd_R87_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, Sw04_command => cmd_R87_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, S126_state => state_S126, S126_lock => S126_locking, S126_command => cmd_R87_S126, J38_state => state_J38, routeState => routes_o(86));
	route_R88 : route_87 port map(clock => clock, routeRequest => routes_i(87), reset => reset, ne292_command => cmd_R88_ne292, ne292_state => state_ne292, ne292_lock => ne292_locking, ne996_command => cmd_R88_ne996, ne996_state => state_ne996, ne996_lock => ne996_locking, Sw04_command => cmd_R88_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, S129_state => state_S129, S129_lock => S129_locking, S129_command => cmd_R88_S129, J37_state => state_J37, routeState => routes_o(87));
	route_R89 : route_88 port map(clock => clock, routeRequest => routes_i(88), reset => reset, ne297_command => cmd_R89_ne297, ne297_state => state_ne297, ne297_lock => ne297_locking, ne996_command => cmd_R89_ne996, ne996_state => state_ne996, ne996_lock => ne996_locking, ne997_command => cmd_R89_ne997, ne997_state => state_ne997, ne997_lock => ne997_locking, Sw03_command => cmd_R89_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, Sw04_command => cmd_R89_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, S129_state => state_S129, S129_lock => S129_locking, S129_command => cmd_R89_S129, S71_state => state_S71, routeState => routes_o(88));
	processed <= processing;
end Behavioral;