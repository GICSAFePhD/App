--  route_66.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity route_66 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne63_state : in nodeStates;
			ne63_lock : in objectLock;
			ne63_command : out routeCommands;
			ne124_state : in nodeStates;
			ne124_lock : in objectLock;
			ne124_command : out routeCommands;
			ne421_state : in nodeStates;
			ne421_lock : in objectLock;
			ne421_command : out routeCommands;
			D18_state : in singleSwitchStates;
			D18_lock : in objectLock;
			D18_command : out routeCommands;
			D19_state : in singleSwitchStates;
			D19_lock : in objectLock;
			D19_command : out routeCommands;
			S95_state : in signalStates;
			S95_lock : in objectLock;
			S95_command : out routeCommands;
			T05_state : in signalStates;
			routeState : out std_logic
		);
	end entity route_66;
architecture Behavioral of route_66 is
	component flipFlop is
		port(
			clock : in std_logic;
			reset : in std_logic;
			Q : out std_logic
		);
	end component flipFlop;
	signal restart : std_logic := '0';
	signal Q : std_logic_vector(27 downto 0) := (others => '0');
	signal routingState : routeStates;
	signal ne63_used , ne124_used , ne421_used : std_logic := '0';
begin
	gen : for i in 0 to 26 generate
		inst: flipFlop port map(Q(i),restart,Q(i+1));
	end generate;
	Q(0) <= clock;

	process(clock)
	begin
		if (clock = '1' and clock'Event) then
		case routingState is
			when WAITING_COMMAND =>
				restart <= '0';
				routeState <= '0';
				if (routeRequest = '1') then
					routingState <= RESERVING_TRACKS;
				end if;
			when RESERVING_TRACKS =>
				if (reset = '1' or (Q(0) = '0' and Q(1) = '0' and Q(2) = '0' and Q(3) = '0' and Q(4) = '0' and Q(5) = '0' and Q(6) = '1' and Q(7) = '1' and Q(8) = '0' and Q(9) = '1' and Q(10) = '1' and Q(11) = '1' and Q(12) = '0' and Q(13) = '0' and Q(14) = '0' and Q(15) = '0' and Q(16) = '0' and Q(17) = '1' and Q(18) = '1' and Q(19) = '0' and Q(20) = '1' and Q(21) = '0' and Q(22) = '0' and Q(23) = '0' and Q(24) = '0' and Q(25) = '1' and Q(26) = '0')) then
					restart <= '1';
					routeState <= '0';
					routingState <= WAITING_COMMAND;
				end if;
				if ((ne63_lock = RELEASED and ne124_lock = RELEASED and ne421_lock = RELEASED) and (ne63_state = FREE and ne124_state = FREE and ne421_state = FREE)) then
					ne63_command <= RESERVE;
					ne124_command <= RESERVE;
					ne421_command <= RESERVE;
					restart <= '0';
				end if;
				if (ne63_lock = RESERVED and ne124_lock = RESERVED and ne421_lock = RESERVED)then
					routingState <= LOCKING_TRACKS;
				end if;
			when LOCKING_TRACKS =>
				if (reset = '1' or (Q(0) = '0' and Q(1) = '0' and Q(2) = '0' and Q(3) = '0' and Q(4) = '0' and Q(5) = '0' and Q(6) = '1' and Q(7) = '1' and Q(8) = '0' and Q(9) = '1' and Q(10) = '1' and Q(11) = '1' and Q(12) = '0' and Q(13) = '0' and Q(14) = '0' and Q(15) = '0' and Q(16) = '0' and Q(17) = '1' and Q(18) = '1' and Q(19) = '0' and Q(20) = '1' and Q(21) = '0' and Q(22) = '0' and Q(23) = '0' and Q(24) = '0' and Q(25) = '1' and Q(26) = '0')) then
					restart <= '1';
					routeState <= '0';
					routingState <= WAITING_COMMAND;
				end if;
				if ((ne63_lock = RESERVED and ne124_lock = RESERVED and ne421_lock = RESERVED) and (ne63_state = FREE and ne124_state = FREE and ne421_state = FREE)) then
					ne63_command <= LOCK;
					ne124_command <= LOCK;
					ne421_command <= LOCK;
					restart <= '0';
				end if;
				if (ne63_lock = LOCKED and ne124_lock = LOCKED and ne421_lock = LOCKED)then
					restart <= '1';
					routingState <= RESERVING_INFRASTRUCTURE;
				end if;
			when RESERVING_INFRASTRUCTURE =>
				if (reset = '1' or (Q(0) = '0' and Q(1) = '0' and Q(2) = '0' and Q(3) = '0' and Q(4) = '0' and Q(5) = '0' and Q(6) = '1' and Q(7) = '1' and Q(8) = '0' and Q(9) = '1' and Q(10) = '1' and Q(11) = '1' and Q(12) = '0' and Q(13) = '0' and Q(14) = '0' and Q(15) = '0' and Q(16) = '0' and Q(17) = '1' and Q(18) = '1' and Q(19) = '0' and Q(20) = '1' and Q(21) = '0' and Q(22) = '0' and Q(23) = '0' and Q(24) = '0' and Q(25) = '1' and Q(26) = '0')) then
					restart <= '1';
					routeState <= '0';
					routingState <= RELEASING_TRACKS;
				end if;
				if (D18_lock = RELEASED and D19_lock = RELEASED) then
					D18_command <= RESERVE;
					D19_command <= RESERVE;
					restart <= '0';
				end if;
				if (D18_lock = RESERVED and D19_lock = RESERVED)then
					routingState <= LOCKING_INFRASTRUCTURE;
				end if;
			when LOCKING_INFRASTRUCTURE =>
				if (reset = '1' or (Q(0) = '0' and Q(1) = '0' and Q(2) = '0' and Q(3) = '0' and Q(4) = '0' and Q(5) = '0' and Q(6) = '1' and Q(7) = '1' and Q(8) = '0' and Q(9) = '1' and Q(10) = '1' and Q(11) = '1' and Q(12) = '0' and Q(13) = '0' and Q(14) = '0' and Q(15) = '0' and Q(16) = '0' and Q(17) = '1' and Q(18) = '1' and Q(19) = '0' and Q(20) = '1' and Q(21) = '0' and Q(22) = '0' and Q(23) = '0' and Q(24) = '0' and Q(25) = '1' and Q(26) = '0')) then
					restart <= '1';
					routeState <= '0';
					routingState <= RELEASING_INFRASTRUCTURE;
				end if;
				if (D18_lock = RELEASED and D19_lock = RELEASED and D18_state = REVERSE and D19_state = REVERSE) then
					D18_command <= LOCK;
					D19_command <= LOCK;
					restart <= '0';
				end if;
				if (D18_lock = LOCKED and D19_lock = LOCKED)then
					routingState <= DRIVING_SIGNAL;
				end if;
			when DRIVING_SIGNAL =>
				if (reset = '1' or (Q(0) = '0' and Q(1) = '0' and Q(2) = '0' and Q(3) = '0' and Q(4) = '0' and Q(5) = '0' and Q(6) = '1' and Q(7) = '1' and Q(8) = '0' and Q(9) = '1' and Q(10) = '1' and Q(11) = '1' and Q(12) = '0' and Q(13) = '0' and Q(14) = '0' and Q(15) = '0' and Q(16) = '0' and Q(17) = '1' and Q(18) = '1' and Q(19) = '0' and Q(20) = '1' and Q(21) = '0' and Q(22) = '0' and Q(23) = '0' and Q(24) = '0' and Q(25) = '1' and Q(26) = '0')) then
					restart <= '1';
					routeState <= '0';
					routingState <= RELEASING_INFRASTRUCTURE;
				end if;
				if (S95_lock = RELEASED) then
					S95_command <= RESERVE;
				end if;
				if (S95_lock = RESERVED and S95_state /= RED) then
					restart <= '0';
					routeState <= '1';
					S95_command <= LOCK;
					routingState <= SEQUENTIAL_RELEASE;
				end if;
			when SEQUENTIAL_RELEASE =>
				--- Sequential release
				if (ne63_used = '0' and ne63_state = OCCUPIED) then 
					ne63_used <= '1';
				end if;
				if (ne63_used = '1' and ne63_state = FREE) then
					ne63_used <= '0';
					ne63_command <= RELEASE;
				end if;
				if (ne124_used = '0' and ne124_state = OCCUPIED) then 
					ne124_used <= '1';
				end if;
				if (ne124_used = '1' and ne124_state = FREE) then
					ne124_used <= '0';
					ne124_command <= RELEASE;
				end if;
				if (ne421_used = '0' and ne421_state = OCCUPIED) then 
					ne421_used <= '1';
					--- Finish -> Release all
					routingState <= RELEASING_INFRASTRUCTURE;
				end if;
			when RELEASING_INFRASTRUCTURE =>
				D18_command <= RELEASE;
				D19_command <= RELEASE;
				routeState <= '0';
				routingState <= RELEASING_TRACKS;
			when RELEASING_TRACKS =>
				ne63_command <= RELEASE;
				ne124_command <= RELEASE;
				ne421_command <= RELEASE;
				routeState <= '0';
				routingState <= WAITING_COMMAND;
			when others =>
				routeState <= '0';
				routingState <= WAITING_COMMAND;
		end case;
		end if;
	end process;
end Behavioral;