--  route_33.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity route_33 is
		port(
			clock : in std_logic;
			routeRequest : in std_logic;
			ne96_state : in nodeStates;
			ne96_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_command : out routeCommands;
			routeState : out std_logic
		);
	end entity route_33;
architecture Behavioral of route_33 is
begin
	routeState <= '0';
end Behavioral;