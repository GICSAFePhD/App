--  node_0.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity node_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R1_command : in routeCommands;
			R8_command : in routeCommands;
			R10_command : in routeCommands;
			R13_command : in routeCommands;
			R14_command : in routeCommands;
			R19_command : in routeCommands;
			R23_command : in routeCommands;
			R24_command : in routeCommands;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end entity node_0;
architecture Behavioral of node_0 is
	signal commandState : routeCommands;
begin

	process(clock)
	begin
		if (clock = '1' and clock'Event) then
			if (reset = '1') then
				commandState <= RELEASE;
			else
				if (R1_command = RELEASE and R8_command = RELEASE and R10_command = RELEASE and R13_command = RELEASE and R14_command = RELEASE and R19_command = RELEASE and R23_command = RELEASE and R24_command = RELEASE and R25_command = RELEASE and R26_command = RELEASE) then
					commandState <= RELEASE;
				else
					if (R1_command = RESERVE or R8_command = RESERVE or R10_command = RESERVE or R13_command = RESERVE or R14_command = RESERVE or R19_command = RESERVE or R23_command = RESERVE or R24_command = RESERVE or R25_command = RESERVE or R26_command = RESERVE) then
						commandState <= RESERVE;
					end if;
					if (R1_command = LOCK or R8_command = LOCK or R10_command = LOCK or R13_command = LOCK or R14_command = LOCK or R19_command = LOCK or R23_command = LOCK or R24_command = LOCK or R25_command = LOCK or R26_command = LOCK) then
						commandState <= LOCK;
					end if;
				end if;
			end if;
		end if;
	end process;

	process(commandState)
	begin
		case commandState is
			when RELEASE => -- AUTOMATIC
				locking <= RELEASED;
			when RESERVE => -- DONT CHANGE
				locking <= RESERVED;
			when LOCK => -- DONT CHANGE
				locking <= LOCKED;
			when others =>
				locking <= LOCKED;
		end case;
	end process;

	process(clock)
	begin
		if (clock = '1' and clock'Event) then
			if (ocupation = '1') then
				state <= FREE;
			else
				state <= OCCUPIED;
			end if;
		end if;
	end process;
end Behavioral;