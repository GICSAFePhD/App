--  splitter.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity splitter is
		generic(
			N : natural := 248;
			N_SIGNALS : natural := 82;
			N_LEVELCROSSINGS : natural := 1;
			N_SINGLESWITCHES : natural := 14;
			N_DOUBLEWITCHES : natural := 8;
			N_TRACKCIRCUITS : natural := 53
		);
		port(
			clock : in std_logic;
			packet :  in std_logic_vector(N-1 downto 0);
			processing :  in std_logic;
			processed :  out std_logic;
			ocupation :  out std_logic_vector(N_TRACKCIRCUITS-1 downto 0);
			signals :  out signals_type;
			levelCrossings : out std_logic;
			singleSwitches : out std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			doubleSwitches : out dSwitches_type;
			reset : in std_logic
		);
	end entity splitter;
architecture Behavioral of splitter is
	Signal tc_s : std_logic_vector(53-1 downto 0);
	Signal sig_s_i,sig_s_o : signals_type;
	Signal lc_s_i,lc_s_o : std_logic;
	Signal ssw_s_i,ssw_s_o : std_logic_vector(14-1 downto 0);
	Signal dsw_s_i,dsw_s_o : dSwitches_type;
begin
	process(clock,reset)
	begin
		if (clock = '1' and clock'Event) then
			if (reset = '1') then
				ocupation <= "00000000000000000000000000000000000000000000000000000";
				signals.lsb <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000";
				signals.msb <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000";
				levelCrossings <= '0';
				singleSwitches <= "00000000000000";
				doubleSwitches.lsb <= "00000000";
				doubleSwitches.msb <= "00000000";
				processed <= '0';
			else
				processed <= processing;
				if processing = '1' then
					ocupation(0) <= packet(247);
					ocupation(1) <= packet(246);
					ocupation(2) <= packet(245);
					ocupation(3) <= packet(244);
					ocupation(4) <= packet(243);
					ocupation(5) <= packet(242);
					ocupation(6) <= packet(241);
					ocupation(7) <= packet(240);
					ocupation(8) <= packet(239);
					ocupation(9) <= packet(238);
					ocupation(10) <= packet(237);
					ocupation(11) <= packet(236);
					ocupation(12) <= packet(235);
					ocupation(13) <= packet(234);
					ocupation(14) <= packet(233);
					ocupation(15) <= packet(232);
					ocupation(16) <= packet(231);
					ocupation(17) <= packet(230);
					ocupation(18) <= packet(229);
					ocupation(19) <= packet(228);
					ocupation(20) <= packet(227);
					ocupation(21) <= packet(226);
					ocupation(22) <= packet(225);
					ocupation(23) <= packet(224);
					ocupation(24) <= packet(223);
					ocupation(25) <= packet(222);
					ocupation(26) <= packet(221);
					ocupation(27) <= packet(220);
					ocupation(28) <= packet(219);
					ocupation(29) <= packet(218);
					ocupation(30) <= packet(217);
					ocupation(31) <= packet(216);
					ocupation(32) <= packet(215);
					ocupation(33) <= packet(214);
					ocupation(34) <= packet(213);
					ocupation(35) <= packet(212);
					ocupation(36) <= packet(211);
					ocupation(37) <= packet(210);
					ocupation(38) <= packet(209);
					ocupation(39) <= packet(208);
					ocupation(40) <= packet(207);
					ocupation(41) <= packet(206);
					ocupation(42) <= packet(205);
					ocupation(43) <= packet(204);
					ocupation(44) <= packet(203);
					ocupation(45) <= packet(202);
					ocupation(46) <= packet(201);
					ocupation(47) <= packet(200);
					ocupation(48) <= packet(199);
					ocupation(49) <= packet(198);
					ocupation(50) <= packet(197);
					ocupation(51) <= packet(196);
					ocupation(52) <= packet(195);
					signals.msb(0) <= packet(194);
					signals.lsb(0) <= packet(193);
					signals.msb(1) <= packet(192);
					signals.lsb(1) <= packet(191);
					signals.msb(2) <= packet(190);
					signals.lsb(2) <= packet(189);
					signals.msb(3) <= packet(188);
					signals.lsb(3) <= packet(187);
					signals.msb(4) <= packet(186);
					signals.lsb(4) <= packet(185);
					signals.msb(5) <= packet(184);
					signals.lsb(5) <= packet(183);
					signals.msb(6) <= packet(182);
					signals.lsb(6) <= packet(181);
					signals.msb(7) <= packet(180);
					signals.lsb(7) <= packet(179);
					signals.msb(8) <= packet(178);
					signals.lsb(8) <= packet(177);
					signals.msb(9) <= packet(176);
					signals.lsb(9) <= packet(175);
					signals.msb(10) <= packet(174);
					signals.lsb(10) <= packet(173);
					signals.msb(11) <= packet(172);
					signals.lsb(11) <= packet(171);
					signals.msb(12) <= packet(170);
					signals.lsb(12) <= packet(169);
					signals.msb(13) <= packet(168);
					signals.lsb(13) <= packet(167);
					signals.msb(14) <= packet(166);
					signals.lsb(14) <= packet(165);
					signals.msb(15) <= packet(164);
					signals.lsb(15) <= packet(163);
					signals.msb(16) <= packet(162);
					signals.lsb(16) <= packet(161);
					signals.msb(17) <= packet(160);
					signals.lsb(17) <= packet(159);
					signals.msb(18) <= packet(158);
					signals.lsb(18) <= packet(157);
					signals.msb(19) <= packet(156);
					signals.lsb(19) <= packet(155);
					signals.msb(20) <= packet(154);
					signals.lsb(20) <= packet(153);
					signals.msb(21) <= packet(152);
					signals.lsb(21) <= packet(151);
					signals.msb(22) <= packet(150);
					signals.lsb(22) <= packet(149);
					signals.msb(23) <= packet(148);
					signals.lsb(23) <= packet(147);
					signals.msb(24) <= packet(146);
					signals.lsb(24) <= packet(145);
					signals.msb(25) <= packet(144);
					signals.lsb(25) <= packet(143);
					signals.msb(26) <= packet(142);
					signals.lsb(26) <= packet(141);
					signals.msb(27) <= packet(140);
					signals.lsb(27) <= packet(139);
					signals.msb(28) <= packet(138);
					signals.lsb(28) <= packet(137);
					signals.msb(29) <= packet(136);
					signals.lsb(29) <= packet(135);
					signals.msb(30) <= packet(134);
					signals.lsb(30) <= packet(133);
					signals.msb(31) <= packet(132);
					signals.lsb(31) <= packet(131);
					signals.msb(32) <= packet(130);
					signals.lsb(32) <= packet(129);
					signals.msb(33) <= packet(128);
					signals.lsb(33) <= packet(127);
					signals.msb(34) <= packet(126);
					signals.lsb(34) <= packet(125);
					signals.msb(35) <= packet(124);
					signals.lsb(35) <= packet(123);
					signals.msb(36) <= packet(122);
					signals.lsb(36) <= packet(121);
					signals.msb(37) <= packet(120);
					signals.lsb(37) <= packet(119);
					signals.msb(38) <= packet(118);
					signals.lsb(38) <= packet(117);
					signals.msb(39) <= packet(116);
					signals.lsb(39) <= packet(115);
					signals.msb(40) <= packet(114);
					signals.lsb(40) <= packet(113);
					signals.msb(41) <= packet(112);
					signals.lsb(41) <= packet(111);
					signals.msb(42) <= packet(110);
					signals.lsb(42) <= packet(109);
					signals.msb(43) <= packet(108);
					signals.lsb(43) <= packet(107);
					signals.msb(44) <= packet(106);
					signals.lsb(44) <= packet(105);
					signals.msb(45) <= packet(104);
					signals.lsb(45) <= packet(103);
					signals.msb(46) <= packet(102);
					signals.lsb(46) <= packet(101);
					signals.msb(47) <= packet(100);
					signals.lsb(47) <= packet(99);
					signals.msb(48) <= packet(98);
					signals.lsb(48) <= packet(97);
					signals.msb(49) <= packet(96);
					signals.lsb(49) <= packet(95);
					signals.msb(50) <= packet(94);
					signals.lsb(50) <= packet(93);
					signals.msb(51) <= packet(92);
					signals.lsb(51) <= packet(91);
					signals.msb(52) <= packet(90);
					signals.lsb(52) <= packet(89);
					signals.msb(53) <= packet(88);
					signals.lsb(53) <= packet(87);
					signals.msb(54) <= packet(86);
					signals.lsb(54) <= packet(85);
					signals.msb(55) <= packet(84);
					signals.lsb(55) <= packet(83);
					signals.msb(56) <= packet(82);
					signals.lsb(56) <= packet(81);
					signals.msb(57) <= packet(80);
					signals.lsb(57) <= packet(79);
					signals.msb(58) <= packet(78);
					signals.lsb(58) <= packet(77);
					signals.msb(59) <= packet(76);
					signals.lsb(59) <= packet(75);
					signals.msb(60) <= packet(74);
					signals.lsb(60) <= packet(73);
					signals.msb(61) <= packet(72);
					signals.lsb(61) <= packet(71);
					signals.msb(62) <= packet(70);
					signals.lsb(62) <= packet(69);
					signals.msb(63) <= packet(68);
					signals.lsb(63) <= packet(67);
					signals.msb(64) <= packet(66);
					signals.lsb(64) <= packet(65);
					signals.msb(65) <= packet(64);
					signals.lsb(65) <= packet(63);
					signals.msb(66) <= packet(62);
					signals.lsb(66) <= packet(61);
					signals.msb(67) <= packet(60);
					signals.lsb(67) <= packet(59);
					signals.msb(68) <= packet(58);
					signals.lsb(68) <= packet(57);
					signals.msb(69) <= packet(56);
					signals.lsb(69) <= packet(55);
					signals.msb(70) <= packet(54);
					signals.lsb(70) <= packet(53);
					signals.msb(71) <= packet(52);
					signals.lsb(71) <= packet(51);
					signals.msb(72) <= packet(50);
					signals.lsb(72) <= packet(49);
					signals.msb(73) <= packet(48);
					signals.lsb(73) <= packet(47);
					signals.msb(74) <= packet(46);
					signals.lsb(74) <= packet(45);
					signals.msb(75) <= packet(44);
					signals.lsb(75) <= packet(43);
					signals.msb(76) <= packet(42);
					signals.lsb(76) <= packet(41);
					signals.msb(77) <= packet(40);
					signals.lsb(77) <= packet(39);
					signals.msb(78) <= packet(38);
					signals.lsb(78) <= packet(37);
					signals.msb(79) <= packet(36);
					signals.lsb(79) <= packet(35);
					signals.msb(80) <= packet(34);
					signals.lsb(80) <= packet(33);
					signals.msb(81) <= packet(32);
					signals.lsb(81) <= packet(31);
					levelCrossings <= packet(30);
					singleSwitches(0) <= packet(29);
					singleSwitches(1) <= packet(28);
					singleSwitches(2) <= packet(27);
					singleSwitches(3) <= packet(26);
					singleSwitches(4) <= packet(25);
					singleSwitches(5) <= packet(24);
					singleSwitches(6) <= packet(23);
					singleSwitches(7) <= packet(22);
					singleSwitches(8) <= packet(21);
					singleSwitches(9) <= packet(20);
					singleSwitches(10) <= packet(19);
					singleSwitches(11) <= packet(18);
					singleSwitches(12) <= packet(17);
					singleSwitches(13) <= packet(16);
					doubleSwitches.msb(0) <= packet(15);
					doubleSwitches.lsb(0) <= packet(14);
					doubleSwitches.msb(1) <= packet(13);
					doubleSwitches.lsb(1) <= packet(12);
					doubleSwitches.msb(2) <= packet(11);
					doubleSwitches.lsb(2) <= packet(10);
					doubleSwitches.msb(3) <= packet(9);
					doubleSwitches.lsb(3) <= packet(8);
					doubleSwitches.msb(4) <= packet(7);
					doubleSwitches.lsb(4) <= packet(6);
					doubleSwitches.msb(5) <= packet(5);
					doubleSwitches.lsb(5) <= packet(4);
					doubleSwitches.msb(6) <= packet(3);
					doubleSwitches.lsb(6) <= packet(2);
					doubleSwitches.msb(7) <= packet(1);
					doubleSwitches.lsb(7) <= packet(0);
				end if;
			end if;
		end if;
	end process;
end Behavioral;