--  network.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity network is
		generic(
			N : natural := 329;
			N_SIGNALS : natural := 82;
			N_ROUTES : natural := 91;
			N_LEVELCROSSINGS : natural := 1;
			N_SINGLESWITCHES : natural := 15;
			N_DOUBLEWITCHES : natural := 2;
			N_SCISSORCROSSINGS : natural := 1;
			N_TRACKCIRCUITS : natural := 53
		);
		port(
			clock : in std_logic;
			processing : in std_logic;
			processed : out std_logic;
			ocupation : in std_logic_vector(N_TRACKCIRCUITS-1 downto 0);
			signals_i : in signals_type;
			signals_o : out signals_type;
			routes_i : in std_logic_vector(N_ROUTES-1 downto 0);
			routes_o : out std_logic_vector(N_ROUTES-1 downto 0);
			levelCrossings_i : in std_logic;
			levelCrossings_o : out std_logic;
			singleSwitches_i : in std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			singleSwitches_o : out std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			scissorCrossings_i : in std_logic;
			scissorCrossings_o : out std_logic;
			doubleSwitches_i : in dSwitches_type;
			doubleSwitches_o : out dSwitches_type;
			reset : in std_logic
		);
	end entity network;
architecture Behavioral of network is
	component levelCrossing_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation_ne95 : in std_logic;
			ocupation_ne9 : in std_logic;
			ocupation_ne59 : in std_logic;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Lc01 : out levelCrossingStates;
			lock_Lc01 : out objectLock
		);
	end component levelCrossing_0;
	component singleSwitch_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R23_command : in routeCommands;
			R38_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_68W02 : out singleSwitchStates;
			lock_68W02 : out objectLock
		);
	end component singleSwitch_0;
	component singleSwitch_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R41_command : in routeCommands;
			R42_command : in routeCommands;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_69W03 : out singleSwitchStates;
			lock_69W03 : out objectLock
		);
	end component singleSwitch_1;
	component singleSwitch_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R3_command : in routeCommands;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			R45_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_69W04 : out singleSwitchStates;
			lock_69W04 : out objectLock
		);
	end component singleSwitch_2;
	component singleSwitch_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R36_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R89_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw06 : out singleSwitchStates;
			lock_Sw06 : out objectLock
		);
	end component singleSwitch_3;
	component singleSwitch_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R47_command : in routeCommands;
			R48_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_70W01 : out singleSwitchStates;
			lock_70W01 : out objectLock
		);
	end component singleSwitch_4;
	component singleSwitch_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R27_command : in routeCommands;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			R51_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_70W02 : out singleSwitchStates;
			lock_70W02 : out objectLock
		);
	end component singleSwitch_5;
	component singleSwitch_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R52_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R55_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw08 : out singleSwitchStates;
			lock_Sw08 : out objectLock
		);
	end component singleSwitch_6;
	component singleSwitch_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R54_command : in routeCommands;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R59_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw09 : out singleSwitchStates;
			lock_Sw09 : out objectLock
		);
	end component singleSwitch_7;
	component singleSwitch_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R7_command : in routeCommands;
			R8_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw12 : out singleSwitchStates;
			lock_Sw12 : out objectLock
		);
	end component singleSwitch_8;
	component singleSwitch_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R5_command : in routeCommands;
			R67_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R77_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw04 : out singleSwitchStates;
			lock_Sw04 : out objectLock
		);
	end component singleSwitch_9;
	component singleSwitch_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R60_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_71W01 : out singleSwitchStates;
			lock_71W01 : out objectLock
		);
	end component singleSwitch_10;
	component singleSwitch_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			R61_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_71W02 : out singleSwitchStates;
			lock_71W02 : out objectLock
		);
	end component singleSwitch_11;
	component singleSwitch_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw11 : out singleSwitchStates;
			lock_Sw11 : out objectLock
		);
	end component singleSwitch_12;
	component singleSwitch_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R8_command : in routeCommands;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw13 : out singleSwitchStates;
			lock_Sw13 : out objectLock
		);
	end component singleSwitch_13;
	component singleSwitch_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R6_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw41 : out singleSwitchStates;
			lock_Sw41 : out objectLock
		);
	end component singleSwitch_14;
	component scissorCrossing_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R14_command : in routeCommands;
			R81_command : in routeCommands;
			R88_command : in routeCommands;
			R91_command : in routeCommands;
			indication : in std_logic;
			command : out std_logic;
			correspondence_Sw03 : out scissorCrossingStates;
			lock_Sw03 : out objectLock
		);
	end component scissorCrossing_0;
	component doubleSwitch_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R5_command : in routeCommands;
			R6_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			indication : in dSwitch_type;
			command : out dSwitch_type;
			correspondence_Sw05 : out doubleSwitchStates;
			lock_Sw05 : out objectLock
		);
	end component doubleSwitch_0;
	component doubleSwitch_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R36_command : in routeCommands;
			R37_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			R89_command : in routeCommands;
			R90_command : in routeCommands;
			indication : in dSwitch_type;
			command : out dSwitch_type;
			correspondence_Sw07 : out doubleSwitchStates;
			lock_Sw07 : out objectLock
		);
	end component doubleSwitch_1;
	component railwaySignal_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne1 : in std_logic;
			correspondence_T01 : out signalStates;
			lock_T01 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_0;
	component railwaySignal_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R1_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne1 : in std_logic;
			correspondence_T02 : out signalStates;
			lock_T02 : out objectLock;
			correspondence_C78 : in signalStates;
			--Ocupation level 2
			ocupation_ne9 : in std_logic;
			correspondence_J46 : in signalStates;
			s68W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_1;
	component railwaySignal_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R38_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne1 : in std_logic;
			correspondence_C78 : out signalStates;
			lock_C78 : out objectLock;
			--Ocupation level 1
			ocupation_ne9 : in std_logic;
			correspondence_J46 : in signalStates;
			s68W02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne95 : in std_logic;
			correspondence_L35 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_2;
	component railwaySignal_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne4 : in std_logic;
			correspondence_T03 : out signalStates;
			lock_T03 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_3;
	component railwaySignal_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R10_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne4 : in std_logic;
			correspondence_L25 : out signalStates;
			lock_L25 : out objectLock;
			--Ocupation level 1
			ocupation_ne106 : in std_logic;
			correspondence_L42 : in signalStates;
			--Ocupation level 2
			ocupation_ne99 : in std_logic;
			correspondence_P68 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_4;
	component railwaySignal_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne7 : in std_logic;
			correspondence_T05 : out signalStates;
			lock_T05 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_5;
	component railwaySignal_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R2_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne7 : in std_logic;
			correspondence_T06 : out signalStates;
			lock_T06 : out objectLock;
			correspondence_J43 : in signalStates;
			--Ocupation level 2
			ocupation_ne9 : in std_logic;
			correspondence_J46 : in signalStates;
			s68W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_6;
	component railwaySignal_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R23_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne7 : in std_logic;
			correspondence_J43 : out signalStates;
			lock_J43 : out objectLock;
			--Ocupation level 1
			ocupation_ne9 : in std_logic;
			correspondence_J46 : in signalStates;
			s68W02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne95 : in std_logic;
			correspondence_L35 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_7;
	component railwaySignal_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R24_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne9 : in std_logic;
			correspondence_J46 : out signalStates;
			lock_J46 : out objectLock;
			--Ocupation level 1
			ocupation_ne95 : in std_logic;
			correspondence_L35 : in signalStates;
			correspondence_X50 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_8;
	component railwaySignal_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne9 : in std_logic;
			correspondence_S80 : out signalStates;
			lock_S80 : out objectLock;
			--Ocupation level 1
			ocupation_ne1 : in std_logic;
			ocupation_ne7 : in std_logic;
			correspondence_T01 : in signalStates;
			correspondence_T05 : in signalStates;
			s68W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_9;
	component railwaySignal_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne14 : in std_logic;
			correspondence_T07 : out signalStates;
			lock_T07 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_10;
	component railwaySignal_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R3_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne14 : in std_logic;
			correspondence_T08 : out signalStates;
			lock_T08 : out objectLock;
			--Ocupation level 1
			ocupation_ne52 : in std_logic;
			correspondence_S146 : in signalStates;
			s69W04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne77 : in std_logic;
			correspondence_B145 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_11;
	component railwaySignal_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R41_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne17 : in std_logic;
			correspondence_C82 : out signalStates;
			lock_C82 : out objectLock;
			--Ocupation level 1
			ocupation_ne59 : in std_logic;
			ocupation_ne95 : in std_logic;
			correspondence_X51 : in signalStates;
			s69W03_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne9 : in std_logic;
			correspondence_S80 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_12;
	component railwaySignal_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R63_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne17 : in std_logic;
			correspondence_C109 : out signalStates;
			lock_C109 : out objectLock;
			--Ocupation level 1
			ocupation_ne78 : in std_logic;
			correspondence_L33 : in signalStates;
			Sw06_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne93 : in std_logic;
			correspondence_L34 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_13;
	component railwaySignal_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R27_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne23 : in std_logic;
			correspondence_P60 : out signalStates;
			lock_P60 : out objectLock;
			--Ocupation level 1
			ocupation_ne26 : in std_logic;
			correspondence_L27 : in signalStates;
			s70W02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne65 : in std_logic;
			correspondence_L30 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_14;
	component railwaySignal_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R46_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne23 : in std_logic;
			correspondence_B89 : out signalStates;
			lock_B89 : out objectLock;
			--Ocupation level 1
			ocupation_ne64 : in std_logic;
			ocupation_ne103 : in std_logic;
			ocupation_ne67 : in std_logic;
			correspondence_P64 : in signalStates;
			--Ocupation level 2
			ocupation_ne70 : in std_logic;
			correspondence_L32 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_15;
	component railwaySignal_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R28_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne24 : in std_logic;
			correspondence_P63 : out signalStates;
			lock_P63 : out objectLock;
			--Ocupation level 1
			ocupation_ne64 : in std_logic;
			ocupation_ne103 : in std_logic;
			ocupation_ne67 : in std_logic;
			correspondence_P64 : in signalStates;
			--Ocupation level 2
			ocupation_ne70 : in std_logic;
			correspondence_L32 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_16;
	component railwaySignal_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R49_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne24 : in std_logic;
			correspondence_B92 : out signalStates;
			lock_B92 : out objectLock;
			--Ocupation level 1
			ocupation_ne26 : in std_logic;
			correspondence_L27 : in signalStates;
			s70W02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne65 : in std_logic;
			correspondence_L30 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_17;
	component railwaySignal_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R11_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne26 : in std_logic;
			correspondence_L27 : out signalStates;
			lock_L27 : out objectLock;
			--Ocupation level 1
			ocupation_ne65 : in std_logic;
			correspondence_L30 : in signalStates;
			--Ocupation level 2
			ocupation_ne102 : in std_logic;
			correspondence_C104 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_18;
	component railwaySignal_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R50_command : in routeCommands;
			R51_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne26 : in std_logic;
			correspondence_S93 : out signalStates;
			lock_S93 : out objectLock;
			--Ocupation level 1
			ocupation_ne23 : in std_logic;
			ocupation_ne24 : in std_logic;
			correspondence_B89 : in signalStates;
			correspondence_P63 : in signalStates;
			s70W02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne67 : in std_logic;
			ocupation_ne103 : in std_logic;
			ocupation_ne64 : in std_logic;
			correspondence_P64 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_19;
	component railwaySignal_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R53_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne29 : in std_logic;
			correspondence_B96 : out signalStates;
			lock_B96 : out objectLock;
			--Ocupation level 1
			ocupation_ne30 : in std_logic;
			correspondence_S122 : in signalStates;
			Sw08_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne90 : in std_logic;
			ocupation_ne91 : in std_logic;
			ocupation_ne86 : in std_logic;
			ocupation_ne87 : in std_logic;
			ocupation_ne89 : in std_logic;
			correspondence_T19 : in signalStates;
			correspondence_T15 : in signalStates;
			correspondence_T21 : in signalStates;
			Sw12_state : in singleSwitchStates;
			Sw11_state : in singleSwitchStates;
			Sw13_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_20;
	component railwaySignal_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R57_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne29 : in std_logic;
			correspondence_B101 : out signalStates;
			lock_B101 : out objectLock;
			correspondence_B96 : in signalStates;
			--Ocupation level 2
			ocupation_ne30 : in std_logic;
			correspondence_S122 : in signalStates;
			Sw08_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_21;
	component railwaySignal_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R54_command : in routeCommands;
			R55_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne30 : in std_logic;
			correspondence_S97 : out signalStates;
			lock_S97 : out objectLock;
			--Ocupation level 1
			ocupation_ne29 : in std_logic;
			ocupation_ne110 : in std_logic;
			ocupation_ne83 : in std_logic;
			correspondence_C138 : in signalStates;
			correspondence_C114 : in signalStates;
			Sw08_state : in singleSwitchStates;
			Sw09_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne101 : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne44 : in std_logic;
			ocupation_ne32 : in std_logic;
			correspondence_S105 : in signalStates;
			correspondence_C100 : in signalStates;
			Sw41_state : in singleSwitchStates;
			Sw04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_22;
	component railwaySignal_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne30 : in std_logic;
			correspondence_S122 : out signalStates;
			lock_S122 : out objectLock;
			--Ocupation level 1
			ocupation_ne89 : in std_logic;
			ocupation_ne91 : in std_logic;
			ocupation_ne87 : in std_logic;
			ocupation_ne86 : in std_logic;
			ocupation_ne90 : in std_logic;
			correspondence_T19 : in signalStates;
			correspondence_T15 : in signalStates;
			correspondence_T21 : in signalStates;
			Sw12_state : in singleSwitchStates;
			Sw11_state : in singleSwitchStates;
			Sw13_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_23;
	component railwaySignal_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R56_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne32 : in std_logic;
			correspondence_C100 : out signalStates;
			lock_C100 : out objectLock;
			--Ocupation level 1
			ocupation_ne110 : in std_logic;
			correspondence_C138 : in signalStates;
			Sw09_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne101 : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne44 : in std_logic;
			correspondence_S105 : in signalStates;
			Sw41_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_24;
	component railwaySignal_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne32 : in std_logic;
			correspondence_S115 : out signalStates;
			lock_S115 : out objectLock;
			--Ocupation level 1
			ocupation_ne83 : in std_logic;
			ocupation_ne82 : in std_logic;
			ocupation_ne41 : in std_logic;
			ocupation_ne84 : in std_logic;
			correspondence_C95 : in signalStates;
			correspondence_P58 : in signalStates;
			correspondence_T13 : in signalStates;
			Sw04_state : in singleSwitchStates;
			Sw05_state : in doubleSwitchStates;
			--Ocupation level 2
			ocupation_ne30 : in std_logic;
			correspondence_S122 : in signalStates;
			Sw08_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_25;
	component railwaySignal_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne41 : in std_logic;
			correspondence_P58 : out signalStates;
			lock_P58 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_26;
	component railwaySignal_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne41 : in std_logic;
			correspondence_B130 : out signalStates;
			lock_B130 : out objectLock;
			--Ocupation level 1
			ocupation_ne82 : in std_logic;
			ocupation_ne32 : in std_logic;
			ocupation_ne85 : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne101 : in std_logic;
			ocupation_ne44 : in std_logic;
			correspondence_C100 : in signalStates;
			correspondence_S105 : in signalStates;
			Sw04_state : in singleSwitchStates;
			Sw05_state : in doubleSwitchStates;
			Sw41_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne110 : in std_logic;
			ocupation_ne26 : in std_logic;
			ocupation_ne65 : in std_logic;
			ocupation_ne48 : in std_logic;
			ocupation_ne43 : in std_logic;
			ocupation_ne102 : in std_logic;
			correspondence_C138 : in signalStates;
			correspondence_L29 : in signalStates;
			correspondence_S93 : in signalStates;
			Sw09_state : in singleSwitchStates;
			s71W01_state : in singleSwitchStates;
			s71W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_27;
	component railwaySignal_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R12_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne44 : in std_logic;
			correspondence_L28 : out signalStates;
			lock_L28 : out objectLock;
			--Ocupation level 1
			ocupation_ne101 : in std_logic;
			correspondence_L40 : in signalStates;
			--Ocupation level 2
			ocupation_ne100 : in std_logic;
			correspondence_S139 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_28;
	component railwaySignal_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne44 : in std_logic;
			correspondence_S105 : out signalStates;
			lock_S105 : out objectLock;
			--Ocupation level 1
			ocupation_ne43 : in std_logic;
			ocupation_ne48 : in std_logic;
			ocupation_ne102 : in std_logic;
			ocupation_ne65 : in std_logic;
			ocupation_ne26 : in std_logic;
			correspondence_L29 : in signalStates;
			correspondence_S93 : in signalStates;
			s71W01_state : in singleSwitchStates;
			s71W02_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne23 : in std_logic;
			ocupation_ne24 : in std_logic;
			correspondence_B89 : in signalStates;
			correspondence_P63 : in signalStates;
			s70W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_29;
	component railwaySignal_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne47 : in std_logic;
			correspondence_T11 : out signalStates;
			lock_T11 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_30;
	component railwaySignal_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne47 : in std_logic;
			correspondence_T12 : out signalStates;
			lock_T12 : out objectLock;
			--Ocupation level 1
			ocupation_ne48 : in std_logic;
			correspondence_L29 : in signalStates;
			s71W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_31;
	component railwaySignal_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne48 : in std_logic;
			correspondence_L29 : out signalStates;
			lock_L29 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_32;
	component railwaySignal_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R42_command : in routeCommands;
			R43_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne59 : in std_logic;
			correspondence_S83 : out signalStates;
			lock_S83 : out objectLock;
			--Ocupation level 1
			ocupation_ne11 : in std_logic;
			ocupation_ne52 : in std_logic;
			ocupation_ne17 : in std_logic;
			correspondence_S146 : in signalStates;
			correspondence_C109 : in signalStates;
			s69W03_state : in singleSwitchStates;
			s69W04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne77 : in std_logic;
			ocupation_ne78 : in std_logic;
			correspondence_B145 : in signalStates;
			correspondence_L33 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			Sw06_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_33;
	component railwaySignal_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R47_command : in routeCommands;
			R48_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne64 : in std_logic;
			correspondence_S90 : out signalStates;
			lock_S90 : out objectLock;
			--Ocupation level 1
			ocupation_ne23 : in std_logic;
			ocupation_ne24 : in std_logic;
			correspondence_P60 : in signalStates;
			correspondence_B92 : in signalStates;
			s70W01_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne26 : in std_logic;
			correspondence_L27 : in signalStates;
			s70W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_34;
	component railwaySignal_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R13_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne65 : in std_logic;
			correspondence_L30 : out signalStates;
			lock_L30 : out objectLock;
			--Ocupation level 1
			ocupation_ne102 : in std_logic;
			correspondence_C104 : in signalStates;
			--Ocupation level 2
			ocupation_ne44 : in std_logic;
			correspondence_L28 : in signalStates;
			s71W01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_35;
	component railwaySignal_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R29_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne67 : in std_logic;
			correspondence_P64 : out signalStates;
			lock_P64 : out objectLock;
			--Ocupation level 1
			ocupation_ne70 : in std_logic;
			correspondence_L32 : in signalStates;
			--Ocupation level 2
			ocupation_ne104 : in std_logic;
			ocupation_ne21 : in std_logic;
			correspondence_P73 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_36;
	component railwaySignal_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R30_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne67 : in std_logic;
			correspondence_P65 : out signalStates;
			lock_P65 : out objectLock;
			--Ocupation level 1
			ocupation_ne103 : in std_logic;
			correspondence_L41 : in signalStates;
			--Ocupation level 2
			ocupation_ne64 : in std_logic;
			correspondence_S90 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_37;
	component railwaySignal_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R14_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne70 : in std_logic;
			correspondence_L32 : out signalStates;
			lock_L32 : out objectLock;
			--Ocupation level 1
			ocupation_ne104 : in std_logic;
			ocupation_ne21 : in std_logic;
			correspondence_P73 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			--Ocupation level 2
			ocupation_ne94 : in std_logic;
			ocupation_ne79 : in std_logic;
			ocupation_ne78 : in std_logic;
			ocupation_ne99 : in std_logic;
			ocupation_ne97 : in std_logic;
			correspondence_L33 : in signalStates;
			correspondence_P69 : in signalStates;
			Sw06_state : in singleSwitchStates;
			Sw07_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_38;
	component railwaySignal_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R15_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne78 : in std_logic;
			correspondence_L33 : out signalStates;
			lock_L33 : out objectLock;
			--Ocupation level 1
			ocupation_ne93 : in std_logic;
			correspondence_L34 : in signalStates;
			--Ocupation level 2
			ocupation_ne96 : in std_logic;
			correspondence_P71 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_39;
	component railwaySignal_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R64_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne78 : in std_logic;
			correspondence_S110 : out signalStates;
			lock_S110 : out objectLock;
			--Ocupation level 1
			ocupation_ne17 : in std_logic;
			ocupation_ne79 : in std_logic;
			ocupation_ne77 : in std_logic;
			ocupation_ne21 : in std_logic;
			correspondence_C82 : in signalStates;
			correspondence_B133 : in signalStates;
			correspondence_P72 : in signalStates;
			Sw06_state : in singleSwitchStates;
			Sw07_state : in doubleSwitchStates;
			--Ocupation level 2
			ocupation_ne95 : in std_logic;
			ocupation_ne59 : in std_logic;
			ocupation_ne52 : in std_logic;
			correspondence_X51 : in signalStates;
			correspondence_S86 : in signalStates;
			correspondence_S144 : in signalStates;
			s69W03_state : in singleSwitchStates;
			Sw03_state : in scissorCrossingStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_40;
	component railwaySignal_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R52_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne83 : in std_logic;
			correspondence_C95 : out signalStates;
			lock_C95 : out objectLock;
			--Ocupation level 1
			ocupation_ne30 : in std_logic;
			correspondence_S122 : in signalStates;
			Sw08_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne90 : in std_logic;
			ocupation_ne91 : in std_logic;
			ocupation_ne86 : in std_logic;
			ocupation_ne87 : in std_logic;
			ocupation_ne89 : in std_logic;
			correspondence_T19 : in signalStates;
			correspondence_T15 : in signalStates;
			correspondence_T21 : in signalStates;
			Sw12_state : in singleSwitchStates;
			Sw11_state : in singleSwitchStates;
			Sw13_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_41;
	component railwaySignal_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R67_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne83 : in std_logic;
			correspondence_C114 : out signalStates;
			lock_C114 : out objectLock;
			--Ocupation level 1
			ocupation_ne32 : in std_logic;
			correspondence_C100 : in signalStates;
			Sw04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne110 : in std_logic;
			correspondence_C138 : in signalStates;
			Sw09_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_42;
	component railwaySignal_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne84 : in std_logic;
			correspondence_T13 : out signalStates;
			lock_T13 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_43;
	component railwaySignal_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R5_command : in routeCommands;
			R6_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne84 : in std_logic;
			correspondence_T14 : out signalStates;
			lock_T14 : out objectLock;
			--Ocupation level 1
			ocupation_ne82 : in std_logic;
			ocupation_ne32 : in std_logic;
			ocupation_ne85 : in std_logic;
			ocupation_ne100 : in std_logic;
			ocupation_ne101 : in std_logic;
			ocupation_ne44 : in std_logic;
			correspondence_C100 : in signalStates;
			correspondence_S105 : in signalStates;
			Sw04_state : in singleSwitchStates;
			Sw05_state : in doubleSwitchStates;
			Sw41_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne110 : in std_logic;
			ocupation_ne26 : in std_logic;
			ocupation_ne65 : in std_logic;
			ocupation_ne48 : in std_logic;
			ocupation_ne43 : in std_logic;
			ocupation_ne102 : in std_logic;
			correspondence_C138 : in signalStates;
			correspondence_L29 : in signalStates;
			correspondence_S93 : in signalStates;
			Sw09_state : in singleSwitchStates;
			s71W01_state : in singleSwitchStates;
			s71W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_44;
	component railwaySignal_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne86 : in std_logic;
			correspondence_T15 : out signalStates;
			lock_T15 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_45;
	component railwaySignal_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R72_command : in routeCommands;
			R73_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne86 : in std_logic;
			correspondence_S119 : out signalStates;
			lock_S119 : out objectLock;
			--Ocupation level 1
			ocupation_ne88 : in std_logic;
			ocupation_ne87 : in std_logic;
			ocupation_ne91 : in std_logic;
			ocupation_ne30 : in std_logic;
			correspondence_T17 : in signalStates;
			correspondence_S97 : in signalStates;
			Sw11_state : in singleSwitchStates;
			Sw12_state : in singleSwitchStates;
			Sw13_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne29 : in std_logic;
			ocupation_ne110 : in std_logic;
			ocupation_ne83 : in std_logic;
			correspondence_C138 : in signalStates;
			correspondence_C114 : in signalStates;
			Sw08_state : in singleSwitchStates;
			Sw09_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_46;
	component railwaySignal_47 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne88 : in std_logic;
			correspondence_T17 : out signalStates;
			lock_T17 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_47;
	component railwaySignal_48 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R71_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne88 : in std_logic;
			correspondence_C118 : out signalStates;
			lock_C118 : out objectLock;
			--Ocupation level 1
			ocupation_ne86 : in std_logic;
			correspondence_T15 : in signalStates;
			Sw11_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_48;
	component railwaySignal_49 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne89 : in std_logic;
			correspondence_T19 : out signalStates;
			lock_T19 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_49;
	component railwaySignal_50 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R7_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne89 : in std_logic;
			correspondence_T20 : out signalStates;
			lock_T20 : out objectLock;
			--Ocupation level 1
			ocupation_ne30 : in std_logic;
			correspondence_S97 : in signalStates;
			Sw12_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne29 : in std_logic;
			ocupation_ne110 : in std_logic;
			ocupation_ne83 : in std_logic;
			correspondence_C138 : in signalStates;
			correspondence_C114 : in signalStates;
			Sw08_state : in singleSwitchStates;
			Sw09_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_50;
	component railwaySignal_51 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne90 : in std_logic;
			correspondence_T21 : out signalStates;
			lock_T21 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_51;
	component railwaySignal_52 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R8_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne90 : in std_logic;
			correspondence_T22 : out signalStates;
			lock_T22 : out objectLock;
			--Ocupation level 1
			ocupation_ne91 : in std_logic;
			ocupation_ne30 : in std_logic;
			correspondence_S97 : in signalStates;
			Sw12_state : in singleSwitchStates;
			Sw13_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne29 : in std_logic;
			ocupation_ne110 : in std_logic;
			ocupation_ne83 : in std_logic;
			correspondence_C138 : in signalStates;
			correspondence_C114 : in signalStates;
			Sw08_state : in singleSwitchStates;
			Sw09_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_52;
	component railwaySignal_53 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R16_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne93 : in std_logic;
			correspondence_L34 : out signalStates;
			lock_L34 : out objectLock;
			--Ocupation level 1
			ocupation_ne96 : in std_logic;
			correspondence_P71 : in signalStates;
			--Ocupation level 2
			ocupation_ne98 : in std_logic;
			correspondence_L38 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_53;
	component railwaySignal_54 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne94 : in std_logic;
			correspondence_S135 : out signalStates;
			lock_S135 : out objectLock;
			--Ocupation level 1
			ocupation_ne77 : in std_logic;
			ocupation_ne21 : in std_logic;
			correspondence_B133 : in signalStates;
			correspondence_P72 : in signalStates;
			Sw07_state : in doubleSwitchStates;
			--Ocupation level 2
			ocupation_ne52 : in std_logic;
			correspondence_S86 : in signalStates;
			correspondence_S144 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_54;
	component railwaySignal_55 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R17_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne95 : in std_logic;
			correspondence_L35 : out signalStates;
			lock_L35 : out objectLock;
			correspondence_X50 : in signalStates;
			--Ocupation level 2
			ocupation_ne59 : in std_logic;
			correspondence_S83 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_55;
	component railwaySignal_56 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R25_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne95 : in std_logic;
			correspondence_X50 : out signalStates;
			lock_X50 : out objectLock;
			--Ocupation level 1
			ocupation_ne59 : in std_logic;
			correspondence_S83 : in signalStates;
			--Ocupation level 2
			ocupation_ne11 : in std_logic;
			ocupation_ne17 : in std_logic;
			ocupation_ne52 : in std_logic;
			correspondence_S146 : in signalStates;
			correspondence_C109 : in signalStates;
			s69W03_state : in singleSwitchStates;
			s69W04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_56;
	component railwaySignal_57 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R26_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne95 : in std_logic;
			correspondence_X51 : out signalStates;
			lock_X51 : out objectLock;
			--Ocupation level 1
			ocupation_ne9 : in std_logic;
			correspondence_S80 : in signalStates;
			--Ocupation level 2
			ocupation_ne1 : in std_logic;
			ocupation_ne7 : in std_logic;
			correspondence_T01 : in signalStates;
			correspondence_T05 : in signalStates;
			s68W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_57;
	component railwaySignal_58 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R33_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne96 : in std_logic;
			correspondence_P70 : out signalStates;
			lock_P70 : out objectLock;
			--Ocupation level 1
			ocupation_ne93 : in std_logic;
			ocupation_ne78 : in std_logic;
			correspondence_S110 : in signalStates;
			--Ocupation level 2
			ocupation_ne79 : in std_logic;
			ocupation_ne21 : in std_logic;
			ocupation_ne17 : in std_logic;
			ocupation_ne77 : in std_logic;
			correspondence_C82 : in signalStates;
			correspondence_B133 : in signalStates;
			correspondence_P72 : in signalStates;
			Sw06_state : in singleSwitchStates;
			Sw07_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_58;
	component railwaySignal_59 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R34_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne96 : in std_logic;
			correspondence_P71 : out signalStates;
			lock_P71 : out objectLock;
			--Ocupation level 1
			ocupation_ne98 : in std_logic;
			correspondence_L38 : in signalStates;
			--Ocupation level 2
			ocupation_ne105 : in std_logic;
			correspondence_T23 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_59;
	component railwaySignal_60 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R18_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne97 : in std_logic;
			correspondence_L37 : out signalStates;
			lock_L37 : out objectLock;
			--Ocupation level 1
			ocupation_ne94 : in std_logic;
			correspondence_S135 : in signalStates;
			--Ocupation level 2
			ocupation_ne21 : in std_logic;
			ocupation_ne77 : in std_logic;
			correspondence_B133 : in signalStates;
			correspondence_P72 : in signalStates;
			Sw07_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_60;
	component railwaySignal_61 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R19_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne98 : in std_logic;
			correspondence_L38 : out signalStates;
			lock_L38 : out objectLock;
			--Ocupation level 1
			ocupation_ne105 : in std_logic;
			correspondence_T23 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_61;
	component railwaySignal_62 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R31_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne99 : in std_logic;
			correspondence_P68 : out signalStates;
			lock_P68 : out objectLock;
			--Ocupation level 1
			ocupation_ne97 : in std_logic;
			correspondence_L37 : in signalStates;
			--Ocupation level 2
			ocupation_ne94 : in std_logic;
			correspondence_S135 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_62;
	component railwaySignal_63 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R32_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne99 : in std_logic;
			correspondence_P69 : out signalStates;
			lock_P69 : out objectLock;
			--Ocupation level 1
			ocupation_ne106 : in std_logic;
			ocupation_ne4 : in std_logic;
			correspondence_T03 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_63;
	component railwaySignal_64 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne100 : in std_logic;
			correspondence_S139 : out signalStates;
			lock_S139 : out objectLock;
			--Ocupation level 1
			ocupation_ne110 : in std_logic;
			ocupation_ne85 : in std_logic;
			correspondence_S102 : in signalStates;
			correspondence_S131 : in signalStates;
			Sw41_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne29 : in std_logic;
			ocupation_ne32 : in std_logic;
			ocupation_ne41 : in std_logic;
			ocupation_ne84 : in std_logic;
			correspondence_S115 : in signalStates;
			correspondence_B101 : in signalStates;
			correspondence_P58 : in signalStates;
			correspondence_T13 : in signalStates;
			Sw09_state : in singleSwitchStates;
			Sw05_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_64;
	component railwaySignal_65 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R20_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne101 : in std_logic;
			correspondence_L40 : out signalStates;
			lock_L40 : out objectLock;
			--Ocupation level 1
			ocupation_ne100 : in std_logic;
			correspondence_S139 : in signalStates;
			--Ocupation level 2
			ocupation_ne110 : in std_logic;
			ocupation_ne85 : in std_logic;
			correspondence_S102 : in signalStates;
			correspondence_S131 : in signalStates;
			Sw41_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_65;
	component railwaySignal_66 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R60_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne102 : in std_logic;
			correspondence_C104 : out signalStates;
			lock_C104 : out objectLock;
			--Ocupation level 1
			ocupation_ne44 : in std_logic;
			correspondence_L28 : in signalStates;
			s71W01_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne101 : in std_logic;
			correspondence_L40 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_66;
	component railwaySignal_67 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R21_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne103 : in std_logic;
			correspondence_L41 : out signalStates;
			lock_L41 : out objectLock;
			--Ocupation level 1
			ocupation_ne64 : in std_logic;
			correspondence_S90 : in signalStates;
			--Ocupation level 2
			ocupation_ne23 : in std_logic;
			ocupation_ne24 : in std_logic;
			correspondence_P60 : in signalStates;
			correspondence_B92 : in signalStates;
			s70W01_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_67;
	component railwaySignal_68 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			ocupation_ne105 : in std_logic;
			correspondence_T23 : out signalStates;
			lock_T23 : out objectLock;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_68;
	component railwaySignal_69 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R9_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne105 : in std_logic;
			correspondence_T24 : out signalStates;
			lock_T24 : out objectLock;
			--Ocupation level 1
			ocupation_ne98 : in std_logic;
			ocupation_ne96 : in std_logic;
			correspondence_P70 : in signalStates;
			--Ocupation level 2
			ocupation_ne78 : in std_logic;
			ocupation_ne93 : in std_logic;
			correspondence_S110 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_69;
	component railwaySignal_70 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R22_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne106 : in std_logic;
			correspondence_L42 : out signalStates;
			lock_L42 : out objectLock;
			--Ocupation level 1
			ocupation_ne99 : in std_logic;
			correspondence_P68 : in signalStates;
			--Ocupation level 2
			ocupation_ne97 : in std_logic;
			correspondence_L37 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_70;
	component railwaySignal_71 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne85 : in std_logic;
			correspondence_S131 : out signalStates;
			lock_S131 : out objectLock;
			--Ocupation level 1
			ocupation_ne41 : in std_logic;
			ocupation_ne84 : in std_logic;
			correspondence_P58 : in signalStates;
			correspondence_T13 : in signalStates;
			Sw05_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_71;
	component railwaySignal_72 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R81_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne77 : in std_logic;
			correspondence_B133 : out signalStates;
			lock_B133 : out objectLock;
			--Ocupation level 1
			ocupation_ne52 : in std_logic;
			correspondence_S86 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			--Ocupation level 2
			ocupation_ne95 : in std_logic;
			ocupation_ne11 : in std_logic;
			ocupation_ne14 : in std_logic;
			ocupation_ne59 : in std_logic;
			correspondence_X51 : in signalStates;
			correspondence_T07 : in signalStates;
			s69W03_state : in singleSwitchStates;
			s69W04_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_72;
	component railwaySignal_73 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R89_command : in routeCommands;
			R90_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne77 : in std_logic;
			correspondence_B145 : out signalStates;
			lock_B145 : out objectLock;
			--Ocupation level 1
			ocupation_ne79 : in std_logic;
			ocupation_ne78 : in std_logic;
			ocupation_ne94 : in std_logic;
			ocupation_ne97 : in std_logic;
			ocupation_ne99 : in std_logic;
			correspondence_L33 : in signalStates;
			correspondence_P69 : in signalStates;
			Sw06_state : in singleSwitchStates;
			Sw07_state : in doubleSwitchStates;
			--Ocupation level 2
			ocupation_ne93 : in std_logic;
			ocupation_ne4 : in std_logic;
			ocupation_ne106 : in std_logic;
			correspondence_L34 : in signalStates;
			correspondence_T03 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_73;
	component railwaySignal_74 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R87_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne104 : in std_logic;
			correspondence_B143 : out signalStates;
			lock_B143 : out objectLock;
			--Ocupation level 1
			ocupation_ne70 : in std_logic;
			correspondence_L32 : in signalStates;
			--Ocupation level 2
			ocupation_ne21 : in std_logic;
			correspondence_P73 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_74;
	component railwaySignal_75 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R44_command : in routeCommands;
			R45_command : in routeCommands;
			Lc01_state : in levelCrossingStates;
			--Ocupation level 0
			ocupation_ne52 : in std_logic;
			correspondence_S86 : out signalStates;
			lock_S86 : out objectLock;
			--Ocupation level 1
			ocupation_ne11 : in std_logic;
			ocupation_ne59 : in std_logic;
			ocupation_ne95 : in std_logic;
			ocupation_ne14 : in std_logic;
			correspondence_X51 : in signalStates;
			correspondence_T07 : in signalStates;
			s69W03_state : in singleSwitchStates;
			s69W04_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne9 : in std_logic;
			correspondence_S80 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_75;
	component railwaySignal_76 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R91_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne52 : in std_logic;
			correspondence_S146 : out signalStates;
			lock_S146 : out objectLock;
			--Ocupation level 1
			ocupation_ne77 : in std_logic;
			correspondence_B145 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			--Ocupation level 2
			ocupation_ne94 : in std_logic;
			ocupation_ne79 : in std_logic;
			ocupation_ne78 : in std_logic;
			ocupation_ne99 : in std_logic;
			ocupation_ne97 : in std_logic;
			correspondence_L33 : in signalStates;
			correspondence_P69 : in signalStates;
			Sw06_state : in singleSwitchStates;
			Sw07_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_76;
	component railwaySignal_77 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R35_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne21 : in std_logic;
			correspondence_P72 : out signalStates;
			lock_P72 : out objectLock;
			correspondence_S144 : in signalStates;
			--Ocupation level 2
			ocupation_ne104 : in std_logic;
			correspondence_B143 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_77;
	component railwaySignal_78 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R36_command : in routeCommands;
			R37_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne21 : in std_logic;
			correspondence_P73 : out signalStates;
			lock_P73 : out objectLock;
			--Ocupation level 1
			ocupation_ne79 : in std_logic;
			ocupation_ne78 : in std_logic;
			ocupation_ne94 : in std_logic;
			ocupation_ne97 : in std_logic;
			ocupation_ne99 : in std_logic;
			correspondence_L33 : in signalStates;
			correspondence_P69 : in signalStates;
			Sw06_state : in singleSwitchStates;
			Sw07_state : in doubleSwitchStates;
			--Ocupation level 2
			ocupation_ne93 : in std_logic;
			ocupation_ne4 : in std_logic;
			ocupation_ne106 : in std_logic;
			correspondence_L34 : in signalStates;
			correspondence_T03 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_78;
	component railwaySignal_79 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R88_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne21 : in std_logic;
			correspondence_S144 : out signalStates;
			lock_S144 : out objectLock;
			--Ocupation level 1
			ocupation_ne104 : in std_logic;
			correspondence_B143 : in signalStates;
			Sw03_state : in scissorCrossingStates;
			--Ocupation level 2
			ocupation_ne70 : in std_logic;
			correspondence_L32 : in signalStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_79;
	component railwaySignal_80 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R58_command : in routeCommands;
			R59_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne110 : in std_logic;
			correspondence_S102 : out signalStates;
			lock_S102 : out objectLock;
			--Ocupation level 1
			ocupation_ne32 : in std_logic;
			ocupation_ne29 : in std_logic;
			correspondence_S115 : in signalStates;
			correspondence_B101 : in signalStates;
			Sw09_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne82 : in std_logic;
			ocupation_ne41 : in std_logic;
			ocupation_ne83 : in std_logic;
			ocupation_ne84 : in std_logic;
			correspondence_C95 : in signalStates;
			correspondence_P58 : in signalStates;
			correspondence_T13 : in signalStates;
			correspondence_B96 : in signalStates;
			Sw04_state : in singleSwitchStates;
			Sw05_state : in doubleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_80;
	component railwaySignal_81 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R84_command : in routeCommands;
			--Ocupation level 0
			ocupation_ne110 : in std_logic;
			correspondence_C138 : out signalStates;
			lock_C138 : out objectLock;
			--Ocupation level 1
			ocupation_ne100 : in std_logic;
			ocupation_ne101 : in std_logic;
			ocupation_ne44 : in std_logic;
			correspondence_S105 : in signalStates;
			Sw41_state : in singleSwitchStates;
			--Ocupation level 2
			ocupation_ne26 : in std_logic;
			ocupation_ne65 : in std_logic;
			ocupation_ne48 : in std_logic;
			ocupation_ne43 : in std_logic;
			ocupation_ne102 : in std_logic;
			correspondence_L29 : in signalStates;
			correspondence_S93 : in signalStates;
			s71W01_state : in singleSwitchStates;
			s71W02_state : in singleSwitchStates;
			indication : in signal_type;
			command : out signal_type
		);
	end component railwaySignal_81;
	component node_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R1_command : in routeCommands;
			R38_command : in routeCommands;
			R39_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_0;
	component node_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R10_command : in routeCommands;
			R32_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_1;
	component node_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R2_command : in routeCommands;
			R23_command : in routeCommands;
			R40_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_2;
	component node_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R23_command : in routeCommands;
			R24_command : in routeCommands;
			R26_command : in routeCommands;
			R38_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_3;
	component node_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_4;
	component node_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R3_command : in routeCommands;
			R45_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_5;
	component node_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_6;
	component node_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R27_command : in routeCommands;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			R50_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_7;
	component node_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R28_command : in routeCommands;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R51_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_8;
	component node_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R27_command : in routeCommands;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			R51_command : in routeCommands;
			R62_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_9;
	component node_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R57_command : in routeCommands;
			R59_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_10;
	component node_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R7_command : in routeCommands;
			R8_command : in routeCommands;
			R52_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R55_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_11;
	component node_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R5_command : in routeCommands;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R67_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R77_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_12;
	component node_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R69_command : in routeCommands;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			R79_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_13;
	component node_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R61_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_14;
	component node_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R12_command : in routeCommands;
			R60_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_15;
	component node_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_16;
	component node_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R4_command : in routeCommands;
			R61_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_17;
	component node_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R25_command : in routeCommands;
			R41_command : in routeCommands;
			R42_command : in routeCommands;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_18;
	component node_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R21_command : in routeCommands;
			R28_command : in routeCommands;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			R48_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_19;
	component node_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R11_command : in routeCommands;
			R13_command : in routeCommands;
			R62_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_20;
	component node_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R28_command : in routeCommands;
			R29_command : in routeCommands;
			R30_command : in routeCommands;
			R46_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_21;
	component node_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R14_command : in routeCommands;
			R29_command : in routeCommands;
			R87_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_22;
	component node_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R15_command : in routeCommands;
			R33_command : in routeCommands;
			R36_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R89_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_23;
	component node_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R36_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R89_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_24;
	component node_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R5_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R77_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_25;
	component node_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R52_command : in routeCommands;
			R55_command : in routeCommands;
			R67_command : in routeCommands;
			R68_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_26;
	component node_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R5_command : in routeCommands;
			R6_command : in routeCommands;
			R70_command : in routeCommands;
			R80_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_27;
	component node_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_28;
	component node_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_29;
	component node_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_30;
	component node_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R7_command : in routeCommands;
			R74_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_31;
	component node_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R76_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_32;
	component node_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R8_command : in routeCommands;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_33;
	component node_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R15_command : in routeCommands;
			R16_command : in routeCommands;
			R33_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_34;
	component node_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R18_command : in routeCommands;
			R37_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			R90_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_35;
	component node_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R17_command : in routeCommands;
			R24_command : in routeCommands;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			R41_command : in routeCommands;
			R44_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_36;
	component node_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R9_command : in routeCommands;
			R16_command : in routeCommands;
			R33_command : in routeCommands;
			R34_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_37;
	component node_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R18_command : in routeCommands;
			R31_command : in routeCommands;
			R37_command : in routeCommands;
			R90_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_38;
	component node_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R9_command : in routeCommands;
			R19_command : in routeCommands;
			R34_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_39;
	component node_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R22_command : in routeCommands;
			R31_command : in routeCommands;
			R32_command : in routeCommands;
			R37_command : in routeCommands;
			R90_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_40;
	component node_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R20_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_41;
	component node_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R12_command : in routeCommands;
			R20_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_42;
	component node_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R13_command : in routeCommands;
			R60_command : in routeCommands;
			R62_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_43;
	component node_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R21_command : in routeCommands;
			R28_command : in routeCommands;
			R30_command : in routeCommands;
			R46_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_44;
	component node_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R9_command : in routeCommands;
			R19_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_45;
	component node_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R10_command : in routeCommands;
			R22_command : in routeCommands;
			R32_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_46;
	component node_47 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R6_command : in routeCommands;
			R78_command : in routeCommands;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			R86_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_47;
	component node_48 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R65_command : in routeCommands;
			R81_command : in routeCommands;
			R82_command : in routeCommands;
			R89_command : in routeCommands;
			R90_command : in routeCommands;
			R91_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_48;
	component node_49 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R14_command : in routeCommands;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_49;
	component node_50 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R3_command : in routeCommands;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			R45_command : in routeCommands;
			R81_command : in routeCommands;
			R91_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_50;
	component node_51 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R14_command : in routeCommands;
			R35_command : in routeCommands;
			R36_command : in routeCommands;
			R37_command : in routeCommands;
			R66_command : in routeCommands;
			R83_command : in routeCommands;
			R88_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_51;
	component node_52 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			ocupation : in std_logic;
			R54_command : in routeCommands;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R59_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			state : out nodeStates;
			locking : out objectLock
		);
	end component node_52;
	component route_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne1_state : in nodeStates;
			ne1_lock : in objectLock;
			ne1_command : out routeCommands;
			T02_state : in signalStates;
			T02_lock : in objectLock;
			T02_command : out routeCommands;
			C78_state : in signalStates;
			routeState : out std_logic
		);
	end component route_0;
	component route_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne7_state : in nodeStates;
			ne7_lock : in objectLock;
			ne7_command : out routeCommands;
			T06_state : in signalStates;
			T06_lock : in objectLock;
			T06_command : out routeCommands;
			J43_state : in signalStates;
			routeState : out std_logic
		);
	end component route_1;
	component route_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne14_state : in nodeStates;
			ne14_lock : in objectLock;
			ne14_command : out routeCommands;
			ne52_state : in nodeStates;
			ne52_lock : in objectLock;
			ne52_command : out routeCommands;
			s69W04_state : in singleSwitchStates;
			s69W04_lock : in objectLock;
			s69W04_command : out routeCommands;
			T08_state : in signalStates;
			T08_lock : in objectLock;
			T08_command : out routeCommands;
			S146_state : in signalStates;
			routeState : out std_logic
		);
	end component route_2;
	component route_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne47_state : in nodeStates;
			ne47_lock : in objectLock;
			ne47_command : out routeCommands;
			ne48_state : in nodeStates;
			ne48_lock : in objectLock;
			ne48_command : out routeCommands;
			s71W02_state : in singleSwitchStates;
			s71W02_lock : in objectLock;
			s71W02_command : out routeCommands;
			T12_state : in signalStates;
			T12_lock : in objectLock;
			T12_command : out routeCommands;
			L29_state : in signalStates;
			routeState : out std_logic
		);
	end component route_3;
	component route_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne84_state : in nodeStates;
			ne84_lock : in objectLock;
			ne84_command : out routeCommands;
			ne82_state : in nodeStates;
			ne82_lock : in objectLock;
			ne82_command : out routeCommands;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			T14_state : in signalStates;
			T14_lock : in objectLock;
			T14_command : out routeCommands;
			C100_state : in signalStates;
			routeState : out std_logic
		);
	end component route_4;
	component route_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne84_state : in nodeStates;
			ne84_lock : in objectLock;
			ne84_command : out routeCommands;
			ne85_state : in nodeStates;
			ne85_lock : in objectLock;
			ne85_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			ne44_state : in nodeStates;
			ne44_lock : in objectLock;
			ne44_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			Sw41_state : in singleSwitchStates;
			Sw41_lock : in objectLock;
			Sw41_command : out routeCommands;
			T14_state : in signalStates;
			T14_lock : in objectLock;
			T14_command : out routeCommands;
			S105_state : in signalStates;
			routeState : out std_logic
		);
	end component route_5;
	component route_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne89_state : in nodeStates;
			ne89_lock : in objectLock;
			ne89_command : out routeCommands;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			Sw12_state : in singleSwitchStates;
			Sw12_lock : in objectLock;
			Sw12_command : out routeCommands;
			T20_state : in signalStates;
			T20_lock : in objectLock;
			T20_command : out routeCommands;
			S97_state : in signalStates;
			routeState : out std_logic
		);
	end component route_6;
	component route_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne90_state : in nodeStates;
			ne90_lock : in objectLock;
			ne90_command : out routeCommands;
			ne91_state : in nodeStates;
			ne91_lock : in objectLock;
			ne91_command : out routeCommands;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			Sw12_state : in singleSwitchStates;
			Sw12_lock : in objectLock;
			Sw12_command : out routeCommands;
			Sw13_state : in singleSwitchStates;
			Sw13_lock : in objectLock;
			Sw13_command : out routeCommands;
			T22_state : in signalStates;
			T22_lock : in objectLock;
			T22_command : out routeCommands;
			S97_state : in signalStates;
			routeState : out std_logic
		);
	end component route_7;
	component route_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne105_state : in nodeStates;
			ne105_lock : in objectLock;
			ne105_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			ne96_state : in nodeStates;
			ne96_lock : in objectLock;
			ne96_command : out routeCommands;
			T24_state : in signalStates;
			T24_lock : in objectLock;
			T24_command : out routeCommands;
			P70_state : in signalStates;
			routeState : out std_logic
		);
	end component route_8;
	component route_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne4_state : in nodeStates;
			ne4_lock : in objectLock;
			ne4_command : out routeCommands;
			ne106_state : in nodeStates;
			ne106_lock : in objectLock;
			ne106_command : out routeCommands;
			L25_state : in signalStates;
			L25_lock : in objectLock;
			L25_command : out routeCommands;
			L42_state : in signalStates;
			routeState : out std_logic
		);
	end component route_9;
	component route_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne26_state : in nodeStates;
			ne26_lock : in objectLock;
			ne26_command : out routeCommands;
			ne65_state : in nodeStates;
			ne65_lock : in objectLock;
			ne65_command : out routeCommands;
			L27_state : in signalStates;
			L27_lock : in objectLock;
			L27_command : out routeCommands;
			L30_state : in signalStates;
			routeState : out std_logic
		);
	end component route_10;
	component route_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne44_state : in nodeStates;
			ne44_lock : in objectLock;
			ne44_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			L28_state : in signalStates;
			L28_lock : in objectLock;
			L28_command : out routeCommands;
			L40_state : in signalStates;
			routeState : out std_logic
		);
	end component route_11;
	component route_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne65_state : in nodeStates;
			ne65_lock : in objectLock;
			ne65_command : out routeCommands;
			ne102_state : in nodeStates;
			ne102_lock : in objectLock;
			ne102_command : out routeCommands;
			L30_state : in signalStates;
			L30_lock : in objectLock;
			L30_command : out routeCommands;
			C104_state : in signalStates;
			routeState : out std_logic
		);
	end component route_12;
	component route_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne70_state : in nodeStates;
			ne70_lock : in objectLock;
			ne70_command : out routeCommands;
			ne104_state : in nodeStates;
			ne104_lock : in objectLock;
			ne104_command : out routeCommands;
			ne21_state : in nodeStates;
			ne21_lock : in objectLock;
			ne21_command : out routeCommands;
			Sw03_state : in scissorCrossingStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			L32_state : in signalStates;
			L32_lock : in objectLock;
			L32_command : out routeCommands;
			P73_state : in signalStates;
			routeState : out std_logic
		);
	end component route_13;
	component route_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			ne93_state : in nodeStates;
			ne93_lock : in objectLock;
			ne93_command : out routeCommands;
			L33_state : in signalStates;
			L33_lock : in objectLock;
			L33_command : out routeCommands;
			L34_state : in signalStates;
			routeState : out std_logic
		);
	end component route_14;
	component route_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne93_state : in nodeStates;
			ne93_lock : in objectLock;
			ne93_command : out routeCommands;
			ne96_state : in nodeStates;
			ne96_lock : in objectLock;
			ne96_command : out routeCommands;
			L34_state : in signalStates;
			L34_lock : in objectLock;
			L34_command : out routeCommands;
			P71_state : in signalStates;
			routeState : out std_logic
		);
	end component route_15;
	component route_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne95_state : in nodeStates;
			ne95_lock : in objectLock;
			ne95_command : out routeCommands;
			L35_state : in signalStates;
			L35_lock : in objectLock;
			L35_command : out routeCommands;
			X50_state : in signalStates;
			routeState : out std_logic
		);
	end component route_16;
	component route_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne97_state : in nodeStates;
			ne97_lock : in objectLock;
			ne97_command : out routeCommands;
			ne94_state : in nodeStates;
			ne94_lock : in objectLock;
			ne94_command : out routeCommands;
			L37_state : in signalStates;
			L37_lock : in objectLock;
			L37_command : out routeCommands;
			S135_state : in signalStates;
			routeState : out std_logic
		);
	end component route_17;
	component route_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			ne105_state : in nodeStates;
			ne105_lock : in objectLock;
			ne105_command : out routeCommands;
			L38_state : in signalStates;
			L38_lock : in objectLock;
			L38_command : out routeCommands;
			T23_state : in signalStates;
			routeState : out std_logic
		);
	end component route_18;
	component route_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			L40_state : in signalStates;
			L40_lock : in objectLock;
			L40_command : out routeCommands;
			S139_state : in signalStates;
			routeState : out std_logic
		);
	end component route_19;
	component route_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne103_state : in nodeStates;
			ne103_lock : in objectLock;
			ne103_command : out routeCommands;
			ne64_state : in nodeStates;
			ne64_lock : in objectLock;
			ne64_command : out routeCommands;
			L41_state : in signalStates;
			L41_lock : in objectLock;
			L41_command : out routeCommands;
			S90_state : in signalStates;
			routeState : out std_logic
		);
	end component route_20;
	component route_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne106_state : in nodeStates;
			ne106_lock : in objectLock;
			ne106_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			L42_state : in signalStates;
			L42_lock : in objectLock;
			L42_command : out routeCommands;
			P68_state : in signalStates;
			routeState : out std_logic
		);
	end component route_21;
	component route_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne7_state : in nodeStates;
			ne7_lock : in objectLock;
			ne7_command : out routeCommands;
			ne9_state : in nodeStates;
			ne9_lock : in objectLock;
			ne9_command : out routeCommands;
			s68W02_state : in singleSwitchStates;
			s68W02_lock : in objectLock;
			s68W02_command : out routeCommands;
			J43_state : in signalStates;
			J43_lock : in objectLock;
			J43_command : out routeCommands;
			J46_state : in signalStates;
			routeState : out std_logic
		);
	end component route_22;
	component route_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne9_state : in nodeStates;
			ne9_lock : in objectLock;
			ne9_command : out routeCommands;
			ne95_state : in nodeStates;
			ne95_lock : in objectLock;
			ne95_command : out routeCommands;
			J46_state : in signalStates;
			J46_lock : in objectLock;
			J46_command : out routeCommands;
			L35_state : in signalStates;
			routeState : out std_logic
		);
	end component route_23;
	component route_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne95_state : in nodeStates;
			ne95_lock : in objectLock;
			ne95_command : out routeCommands;
			ne59_state : in nodeStates;
			ne59_lock : in objectLock;
			ne59_command : out routeCommands;
			Lc01_state : in levelCrossingStates;
			Lc01_lock : in objectLock;
			Lc01_command : out routeCommands;
			X50_state : in signalStates;
			X50_lock : in objectLock;
			X50_command : out routeCommands;
			S83_state : in signalStates;
			routeState : out std_logic
		);
	end component route_24;
	component route_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne95_state : in nodeStates;
			ne95_lock : in objectLock;
			ne95_command : out routeCommands;
			ne9_state : in nodeStates;
			ne9_lock : in objectLock;
			ne9_command : out routeCommands;
			Lc01_state : in levelCrossingStates;
			Lc01_lock : in objectLock;
			Lc01_command : out routeCommands;
			X51_state : in signalStates;
			X51_lock : in objectLock;
			X51_command : out routeCommands;
			S80_state : in signalStates;
			routeState : out std_logic
		);
	end component route_25;
	component route_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne23_state : in nodeStates;
			ne23_lock : in objectLock;
			ne23_command : out routeCommands;
			ne26_state : in nodeStates;
			ne26_lock : in objectLock;
			ne26_command : out routeCommands;
			s70W02_state : in singleSwitchStates;
			s70W02_lock : in objectLock;
			s70W02_command : out routeCommands;
			P60_state : in signalStates;
			P60_lock : in objectLock;
			P60_command : out routeCommands;
			L27_state : in signalStates;
			routeState : out std_logic
		);
	end component route_26;
	component route_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne24_state : in nodeStates;
			ne24_lock : in objectLock;
			ne24_command : out routeCommands;
			ne64_state : in nodeStates;
			ne64_lock : in objectLock;
			ne64_command : out routeCommands;
			ne103_state : in nodeStates;
			ne103_lock : in objectLock;
			ne103_command : out routeCommands;
			ne67_state : in nodeStates;
			ne67_lock : in objectLock;
			ne67_command : out routeCommands;
			P63_state : in signalStates;
			P63_lock : in objectLock;
			P63_command : out routeCommands;
			P64_state : in signalStates;
			routeState : out std_logic
		);
	end component route_27;
	component route_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne67_state : in nodeStates;
			ne67_lock : in objectLock;
			ne67_command : out routeCommands;
			ne70_state : in nodeStates;
			ne70_lock : in objectLock;
			ne70_command : out routeCommands;
			P64_state : in signalStates;
			P64_lock : in objectLock;
			P64_command : out routeCommands;
			L32_state : in signalStates;
			routeState : out std_logic
		);
	end component route_28;
	component route_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne67_state : in nodeStates;
			ne67_lock : in objectLock;
			ne67_command : out routeCommands;
			ne103_state : in nodeStates;
			ne103_lock : in objectLock;
			ne103_command : out routeCommands;
			P65_state : in signalStates;
			P65_lock : in objectLock;
			P65_command : out routeCommands;
			L41_state : in signalStates;
			routeState : out std_logic
		);
	end component route_29;
	component route_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			ne97_state : in nodeStates;
			ne97_lock : in objectLock;
			ne97_command : out routeCommands;
			P68_state : in signalStates;
			P68_lock : in objectLock;
			P68_command : out routeCommands;
			L37_state : in signalStates;
			routeState : out std_logic
		);
	end component route_30;
	component route_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			ne106_state : in nodeStates;
			ne106_lock : in objectLock;
			ne106_command : out routeCommands;
			ne4_state : in nodeStates;
			ne4_lock : in objectLock;
			ne4_command : out routeCommands;
			P69_state : in signalStates;
			P69_lock : in objectLock;
			P69_command : out routeCommands;
			T03_state : in signalStates;
			routeState : out std_logic
		);
	end component route_31;
	component route_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne96_state : in nodeStates;
			ne96_lock : in objectLock;
			ne96_command : out routeCommands;
			ne93_state : in nodeStates;
			ne93_lock : in objectLock;
			ne93_command : out routeCommands;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			P70_state : in signalStates;
			P70_lock : in objectLock;
			P70_command : out routeCommands;
			S110_state : in signalStates;
			routeState : out std_logic
		);
	end component route_32;
	component route_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne96_state : in nodeStates;
			ne96_lock : in objectLock;
			ne96_command : out routeCommands;
			ne98_state : in nodeStates;
			ne98_lock : in objectLock;
			ne98_command : out routeCommands;
			P71_state : in signalStates;
			P71_lock : in objectLock;
			P71_command : out routeCommands;
			L38_state : in signalStates;
			routeState : out std_logic
		);
	end component route_33;
	component route_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne21_state : in nodeStates;
			ne21_lock : in objectLock;
			ne21_command : out routeCommands;
			P72_state : in signalStates;
			P72_lock : in objectLock;
			P72_command : out routeCommands;
			S144_state : in signalStates;
			routeState : out std_logic
		);
	end component route_34;
	component route_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne21_state : in nodeStates;
			ne21_lock : in objectLock;
			ne21_command : out routeCommands;
			ne79_state : in nodeStates;
			ne79_lock : in objectLock;
			ne79_command : out routeCommands;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			Sw06_state : in singleSwitchStates;
			Sw06_lock : in objectLock;
			Sw06_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			P73_state : in signalStates;
			P73_lock : in objectLock;
			P73_command : out routeCommands;
			L33_state : in signalStates;
			routeState : out std_logic
		);
	end component route_35;
	component route_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne21_state : in nodeStates;
			ne21_lock : in objectLock;
			ne21_command : out routeCommands;
			ne94_state : in nodeStates;
			ne94_lock : in objectLock;
			ne94_command : out routeCommands;
			ne97_state : in nodeStates;
			ne97_lock : in objectLock;
			ne97_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			P73_state : in signalStates;
			P73_lock : in objectLock;
			P73_command : out routeCommands;
			P69_state : in signalStates;
			routeState : out std_logic
		);
	end component route_36;
	component route_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne1_state : in nodeStates;
			ne1_lock : in objectLock;
			ne1_command : out routeCommands;
			ne9_state : in nodeStates;
			ne9_lock : in objectLock;
			ne9_command : out routeCommands;
			s68W02_state : in singleSwitchStates;
			s68W02_lock : in objectLock;
			s68W02_command : out routeCommands;
			C78_state : in signalStates;
			C78_lock : in objectLock;
			C78_command : out routeCommands;
			J46_state : in signalStates;
			routeState : out std_logic
		);
	end component route_37;
	component route_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne9_state : in nodeStates;
			ne9_lock : in objectLock;
			ne9_command : out routeCommands;
			ne1_state : in nodeStates;
			ne1_lock : in objectLock;
			ne1_command : out routeCommands;
			s68W02_state : in singleSwitchStates;
			s68W02_lock : in objectLock;
			s68W02_command : out routeCommands;
			S80_state : in signalStates;
			S80_lock : in objectLock;
			S80_command : out routeCommands;
			T01_state : in signalStates;
			routeState : out std_logic
		);
	end component route_38;
	component route_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne9_state : in nodeStates;
			ne9_lock : in objectLock;
			ne9_command : out routeCommands;
			ne7_state : in nodeStates;
			ne7_lock : in objectLock;
			ne7_command : out routeCommands;
			s68W02_state : in singleSwitchStates;
			s68W02_lock : in objectLock;
			s68W02_command : out routeCommands;
			S80_state : in signalStates;
			S80_lock : in objectLock;
			S80_command : out routeCommands;
			T05_state : in signalStates;
			routeState : out std_logic
		);
	end component route_39;
	component route_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne17_state : in nodeStates;
			ne17_lock : in objectLock;
			ne17_command : out routeCommands;
			ne59_state : in nodeStates;
			ne59_lock : in objectLock;
			ne59_command : out routeCommands;
			ne95_state : in nodeStates;
			ne95_lock : in objectLock;
			ne95_command : out routeCommands;
			s69W03_state : in singleSwitchStates;
			s69W03_lock : in objectLock;
			s69W03_command : out routeCommands;
			C82_state : in signalStates;
			C82_lock : in objectLock;
			C82_command : out routeCommands;
			X51_state : in signalStates;
			routeState : out std_logic
		);
	end component route_40;
	component route_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne59_state : in nodeStates;
			ne59_lock : in objectLock;
			ne59_command : out routeCommands;
			ne11_state : in nodeStates;
			ne11_lock : in objectLock;
			ne11_command : out routeCommands;
			ne52_state : in nodeStates;
			ne52_lock : in objectLock;
			ne52_command : out routeCommands;
			s69W03_state : in singleSwitchStates;
			s69W03_lock : in objectLock;
			s69W03_command : out routeCommands;
			s69W04_state : in singleSwitchStates;
			s69W04_lock : in objectLock;
			s69W04_command : out routeCommands;
			S83_state : in signalStates;
			S83_lock : in objectLock;
			S83_command : out routeCommands;
			S146_state : in signalStates;
			routeState : out std_logic
		);
	end component route_41;
	component route_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne59_state : in nodeStates;
			ne59_lock : in objectLock;
			ne59_command : out routeCommands;
			ne17_state : in nodeStates;
			ne17_lock : in objectLock;
			ne17_command : out routeCommands;
			s69W03_state : in singleSwitchStates;
			s69W03_lock : in objectLock;
			s69W03_command : out routeCommands;
			S83_state : in signalStates;
			S83_lock : in objectLock;
			S83_command : out routeCommands;
			C109_state : in signalStates;
			routeState : out std_logic
		);
	end component route_42;
	component route_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne52_state : in nodeStates;
			ne52_lock : in objectLock;
			ne52_command : out routeCommands;
			ne11_state : in nodeStates;
			ne11_lock : in objectLock;
			ne11_command : out routeCommands;
			ne59_state : in nodeStates;
			ne59_lock : in objectLock;
			ne59_command : out routeCommands;
			ne95_state : in nodeStates;
			ne95_lock : in objectLock;
			ne95_command : out routeCommands;
			s69W03_state : in singleSwitchStates;
			s69W03_lock : in objectLock;
			s69W03_command : out routeCommands;
			s69W04_state : in singleSwitchStates;
			s69W04_lock : in objectLock;
			s69W04_command : out routeCommands;
			S86_state : in signalStates;
			S86_lock : in objectLock;
			S86_command : out routeCommands;
			X51_state : in signalStates;
			routeState : out std_logic
		);
	end component route_43;
	component route_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne52_state : in nodeStates;
			ne52_lock : in objectLock;
			ne52_command : out routeCommands;
			ne14_state : in nodeStates;
			ne14_lock : in objectLock;
			ne14_command : out routeCommands;
			s69W04_state : in singleSwitchStates;
			s69W04_lock : in objectLock;
			s69W04_command : out routeCommands;
			S86_state : in signalStates;
			S86_lock : in objectLock;
			S86_command : out routeCommands;
			T07_state : in signalStates;
			routeState : out std_logic
		);
	end component route_44;
	component route_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne23_state : in nodeStates;
			ne23_lock : in objectLock;
			ne23_command : out routeCommands;
			ne64_state : in nodeStates;
			ne64_lock : in objectLock;
			ne64_command : out routeCommands;
			ne103_state : in nodeStates;
			ne103_lock : in objectLock;
			ne103_command : out routeCommands;
			ne67_state : in nodeStates;
			ne67_lock : in objectLock;
			ne67_command : out routeCommands;
			B89_state : in signalStates;
			B89_lock : in objectLock;
			B89_command : out routeCommands;
			P64_state : in signalStates;
			routeState : out std_logic
		);
	end component route_45;
	component route_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne64_state : in nodeStates;
			ne64_lock : in objectLock;
			ne64_command : out routeCommands;
			ne23_state : in nodeStates;
			ne23_lock : in objectLock;
			ne23_command : out routeCommands;
			s70W01_state : in singleSwitchStates;
			s70W01_lock : in objectLock;
			s70W01_command : out routeCommands;
			S90_state : in signalStates;
			S90_lock : in objectLock;
			S90_command : out routeCommands;
			P60_state : in signalStates;
			routeState : out std_logic
		);
	end component route_46;
	component route_47 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne64_state : in nodeStates;
			ne64_lock : in objectLock;
			ne64_command : out routeCommands;
			ne24_state : in nodeStates;
			ne24_lock : in objectLock;
			ne24_command : out routeCommands;
			s70W01_state : in singleSwitchStates;
			s70W01_lock : in objectLock;
			s70W01_command : out routeCommands;
			S90_state : in signalStates;
			S90_lock : in objectLock;
			S90_command : out routeCommands;
			B92_state : in signalStates;
			routeState : out std_logic
		);
	end component route_47;
	component route_48 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne24_state : in nodeStates;
			ne24_lock : in objectLock;
			ne24_command : out routeCommands;
			ne26_state : in nodeStates;
			ne26_lock : in objectLock;
			ne26_command : out routeCommands;
			s70W02_state : in singleSwitchStates;
			s70W02_lock : in objectLock;
			s70W02_command : out routeCommands;
			B92_state : in signalStates;
			B92_lock : in objectLock;
			B92_command : out routeCommands;
			L27_state : in signalStates;
			routeState : out std_logic
		);
	end component route_48;
	component route_49 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne26_state : in nodeStates;
			ne26_lock : in objectLock;
			ne26_command : out routeCommands;
			ne23_state : in nodeStates;
			ne23_lock : in objectLock;
			ne23_command : out routeCommands;
			s70W02_state : in singleSwitchStates;
			s70W02_lock : in objectLock;
			s70W02_command : out routeCommands;
			S93_state : in signalStates;
			S93_lock : in objectLock;
			S93_command : out routeCommands;
			B89_state : in signalStates;
			routeState : out std_logic
		);
	end component route_49;
	component route_50 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne26_state : in nodeStates;
			ne26_lock : in objectLock;
			ne26_command : out routeCommands;
			ne24_state : in nodeStates;
			ne24_lock : in objectLock;
			ne24_command : out routeCommands;
			s70W02_state : in singleSwitchStates;
			s70W02_lock : in objectLock;
			s70W02_command : out routeCommands;
			S93_state : in signalStates;
			S93_lock : in objectLock;
			S93_command : out routeCommands;
			P63_state : in signalStates;
			routeState : out std_logic
		);
	end component route_50;
	component route_51 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne83_state : in nodeStates;
			ne83_lock : in objectLock;
			ne83_command : out routeCommands;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			Sw08_state : in singleSwitchStates;
			Sw08_lock : in objectLock;
			Sw08_command : out routeCommands;
			C95_state : in signalStates;
			C95_lock : in objectLock;
			C95_command : out routeCommands;
			S122_state : in signalStates;
			routeState : out std_logic
		);
	end component route_51;
	component route_52 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne29_state : in nodeStates;
			ne29_lock : in objectLock;
			ne29_command : out routeCommands;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			Sw08_state : in singleSwitchStates;
			Sw08_lock : in objectLock;
			Sw08_command : out routeCommands;
			B96_state : in signalStates;
			B96_lock : in objectLock;
			B96_command : out routeCommands;
			S122_state : in signalStates;
			routeState : out std_logic
		);
	end component route_52;
	component route_53 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			ne29_state : in nodeStates;
			ne29_lock : in objectLock;
			ne29_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			Sw08_state : in singleSwitchStates;
			Sw08_lock : in objectLock;
			Sw08_command : out routeCommands;
			Sw09_state : in singleSwitchStates;
			Sw09_lock : in objectLock;
			Sw09_command : out routeCommands;
			S97_state : in signalStates;
			S97_lock : in objectLock;
			S97_command : out routeCommands;
			C138_state : in signalStates;
			routeState : out std_logic
		);
	end component route_53;
	component route_54 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			ne83_state : in nodeStates;
			ne83_lock : in objectLock;
			ne83_command : out routeCommands;
			Sw08_state : in singleSwitchStates;
			Sw08_lock : in objectLock;
			Sw08_command : out routeCommands;
			S97_state : in signalStates;
			S97_lock : in objectLock;
			S97_command : out routeCommands;
			C114_state : in signalStates;
			routeState : out std_logic
		);
	end component route_54;
	component route_55 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			Sw09_state : in singleSwitchStates;
			Sw09_lock : in objectLock;
			Sw09_command : out routeCommands;
			C100_state : in signalStates;
			C100_lock : in objectLock;
			C100_command : out routeCommands;
			C138_state : in signalStates;
			routeState : out std_logic
		);
	end component route_55;
	component route_56 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne29_state : in nodeStates;
			ne29_lock : in objectLock;
			ne29_command : out routeCommands;
			B101_state : in signalStates;
			B101_lock : in objectLock;
			B101_command : out routeCommands;
			B96_state : in signalStates;
			routeState : out std_logic
		);
	end component route_56;
	component route_57 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			Sw09_state : in singleSwitchStates;
			Sw09_lock : in objectLock;
			Sw09_command : out routeCommands;
			S102_state : in signalStates;
			S102_lock : in objectLock;
			S102_command : out routeCommands;
			S115_state : in signalStates;
			routeState : out std_logic
		);
	end component route_57;
	component route_58 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			ne29_state : in nodeStates;
			ne29_lock : in objectLock;
			ne29_command : out routeCommands;
			Sw09_state : in singleSwitchStates;
			Sw09_lock : in objectLock;
			Sw09_command : out routeCommands;
			S102_state : in signalStates;
			S102_lock : in objectLock;
			S102_command : out routeCommands;
			B101_state : in signalStates;
			routeState : out std_logic
		);
	end component route_58;
	component route_59 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne102_state : in nodeStates;
			ne102_lock : in objectLock;
			ne102_command : out routeCommands;
			ne44_state : in nodeStates;
			ne44_lock : in objectLock;
			ne44_command : out routeCommands;
			s71W01_state : in singleSwitchStates;
			s71W01_lock : in objectLock;
			s71W01_command : out routeCommands;
			C104_state : in signalStates;
			C104_lock : in objectLock;
			C104_command : out routeCommands;
			L28_state : in signalStates;
			routeState : out std_logic
		);
	end component route_59;
	component route_60 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne44_state : in nodeStates;
			ne44_lock : in objectLock;
			ne44_command : out routeCommands;
			ne43_state : in nodeStates;
			ne43_lock : in objectLock;
			ne43_command : out routeCommands;
			ne48_state : in nodeStates;
			ne48_lock : in objectLock;
			ne48_command : out routeCommands;
			s71W01_state : in singleSwitchStates;
			s71W01_lock : in objectLock;
			s71W01_command : out routeCommands;
			s71W02_state : in singleSwitchStates;
			s71W02_lock : in objectLock;
			s71W02_command : out routeCommands;
			S105_state : in signalStates;
			S105_lock : in objectLock;
			S105_command : out routeCommands;
			L29_state : in signalStates;
			routeState : out std_logic
		);
	end component route_60;
	component route_61 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne44_state : in nodeStates;
			ne44_lock : in objectLock;
			ne44_command : out routeCommands;
			ne102_state : in nodeStates;
			ne102_lock : in objectLock;
			ne102_command : out routeCommands;
			ne65_state : in nodeStates;
			ne65_lock : in objectLock;
			ne65_command : out routeCommands;
			ne26_state : in nodeStates;
			ne26_lock : in objectLock;
			ne26_command : out routeCommands;
			s71W01_state : in singleSwitchStates;
			s71W01_lock : in objectLock;
			s71W01_command : out routeCommands;
			S105_state : in signalStates;
			S105_lock : in objectLock;
			S105_command : out routeCommands;
			S93_state : in signalStates;
			routeState : out std_logic
		);
	end component route_61;
	component route_62 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne17_state : in nodeStates;
			ne17_lock : in objectLock;
			ne17_command : out routeCommands;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			Sw06_state : in singleSwitchStates;
			Sw06_lock : in objectLock;
			Sw06_command : out routeCommands;
			C109_state : in signalStates;
			C109_lock : in objectLock;
			C109_command : out routeCommands;
			L33_state : in signalStates;
			routeState : out std_logic
		);
	end component route_62;
	component route_63 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			ne17_state : in nodeStates;
			ne17_lock : in objectLock;
			ne17_command : out routeCommands;
			Sw06_state : in singleSwitchStates;
			Sw06_lock : in objectLock;
			Sw06_command : out routeCommands;
			S110_state : in signalStates;
			S110_lock : in objectLock;
			S110_command : out routeCommands;
			C82_state : in signalStates;
			routeState : out std_logic
		);
	end component route_63;
	component route_64 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			ne79_state : in nodeStates;
			ne79_lock : in objectLock;
			ne79_command : out routeCommands;
			ne77_state : in nodeStates;
			ne77_lock : in objectLock;
			ne77_command : out routeCommands;
			Sw06_state : in singleSwitchStates;
			Sw06_lock : in objectLock;
			Sw06_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			S110_state : in signalStates;
			S110_lock : in objectLock;
			S110_command : out routeCommands;
			B133_state : in signalStates;
			routeState : out std_logic
		);
	end component route_64;
	component route_65 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			ne79_state : in nodeStates;
			ne79_lock : in objectLock;
			ne79_command : out routeCommands;
			ne21_state : in nodeStates;
			ne21_lock : in objectLock;
			ne21_command : out routeCommands;
			Sw06_state : in singleSwitchStates;
			Sw06_lock : in objectLock;
			Sw06_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			S110_state : in signalStates;
			S110_lock : in objectLock;
			S110_command : out routeCommands;
			P72_state : in signalStates;
			routeState : out std_logic
		);
	end component route_65;
	component route_66 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne83_state : in nodeStates;
			ne83_lock : in objectLock;
			ne83_command : out routeCommands;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			C114_state : in signalStates;
			C114_lock : in objectLock;
			C114_command : out routeCommands;
			C100_state : in signalStates;
			routeState : out std_logic
		);
	end component route_66;
	component route_67 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			ne83_state : in nodeStates;
			ne83_lock : in objectLock;
			ne83_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			S115_state : in signalStates;
			S115_lock : in objectLock;
			S115_command : out routeCommands;
			C95_state : in signalStates;
			routeState : out std_logic
		);
	end component route_67;
	component route_68 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			ne82_state : in nodeStates;
			ne82_lock : in objectLock;
			ne82_command : out routeCommands;
			ne41_state : in nodeStates;
			ne41_lock : in objectLock;
			ne41_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			S115_state : in signalStates;
			S115_lock : in objectLock;
			S115_command : out routeCommands;
			P58_state : in signalStates;
			routeState : out std_logic
		);
	end component route_68;
	component route_69 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			ne82_state : in nodeStates;
			ne82_lock : in objectLock;
			ne82_command : out routeCommands;
			ne84_state : in nodeStates;
			ne84_lock : in objectLock;
			ne84_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			S115_state : in signalStates;
			S115_lock : in objectLock;
			S115_command : out routeCommands;
			T13_state : in signalStates;
			routeState : out std_logic
		);
	end component route_69;
	component route_70 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne88_state : in nodeStates;
			ne88_lock : in objectLock;
			ne88_command : out routeCommands;
			ne86_state : in nodeStates;
			ne86_lock : in objectLock;
			ne86_command : out routeCommands;
			Sw11_state : in singleSwitchStates;
			Sw11_lock : in objectLock;
			Sw11_command : out routeCommands;
			C118_state : in signalStates;
			C118_lock : in objectLock;
			C118_command : out routeCommands;
			T15_state : in signalStates;
			routeState : out std_logic
		);
	end component route_70;
	component route_71 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne86_state : in nodeStates;
			ne86_lock : in objectLock;
			ne86_command : out routeCommands;
			ne88_state : in nodeStates;
			ne88_lock : in objectLock;
			ne88_command : out routeCommands;
			Sw11_state : in singleSwitchStates;
			Sw11_lock : in objectLock;
			Sw11_command : out routeCommands;
			S119_state : in signalStates;
			S119_lock : in objectLock;
			S119_command : out routeCommands;
			T17_state : in signalStates;
			routeState : out std_logic
		);
	end component route_71;
	component route_72 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne86_state : in nodeStates;
			ne86_lock : in objectLock;
			ne86_command : out routeCommands;
			ne87_state : in nodeStates;
			ne87_lock : in objectLock;
			ne87_command : out routeCommands;
			ne91_state : in nodeStates;
			ne91_lock : in objectLock;
			ne91_command : out routeCommands;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			Sw11_state : in singleSwitchStates;
			Sw11_lock : in objectLock;
			Sw11_command : out routeCommands;
			Sw12_state : in singleSwitchStates;
			Sw12_lock : in objectLock;
			Sw12_command : out routeCommands;
			Sw13_state : in singleSwitchStates;
			Sw13_lock : in objectLock;
			Sw13_command : out routeCommands;
			S119_state : in signalStates;
			S119_lock : in objectLock;
			S119_command : out routeCommands;
			S97_state : in signalStates;
			routeState : out std_logic
		);
	end component route_72;
	component route_73 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			ne89_state : in nodeStates;
			ne89_lock : in objectLock;
			ne89_command : out routeCommands;
			Sw12_state : in singleSwitchStates;
			Sw12_lock : in objectLock;
			Sw12_command : out routeCommands;
			S122_state : in signalStates;
			S122_lock : in objectLock;
			S122_command : out routeCommands;
			T19_state : in signalStates;
			routeState : out std_logic
		);
	end component route_73;
	component route_74 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			ne91_state : in nodeStates;
			ne91_lock : in objectLock;
			ne91_command : out routeCommands;
			ne87_state : in nodeStates;
			ne87_lock : in objectLock;
			ne87_command : out routeCommands;
			ne86_state : in nodeStates;
			ne86_lock : in objectLock;
			ne86_command : out routeCommands;
			Sw11_state : in singleSwitchStates;
			Sw11_lock : in objectLock;
			Sw11_command : out routeCommands;
			Sw12_state : in singleSwitchStates;
			Sw12_lock : in objectLock;
			Sw12_command : out routeCommands;
			Sw13_state : in singleSwitchStates;
			Sw13_lock : in objectLock;
			Sw13_command : out routeCommands;
			S122_state : in signalStates;
			S122_lock : in objectLock;
			S122_command : out routeCommands;
			T15_state : in signalStates;
			routeState : out std_logic
		);
	end component route_74;
	component route_75 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne30_state : in nodeStates;
			ne30_lock : in objectLock;
			ne30_command : out routeCommands;
			ne91_state : in nodeStates;
			ne91_lock : in objectLock;
			ne91_command : out routeCommands;
			ne90_state : in nodeStates;
			ne90_lock : in objectLock;
			ne90_command : out routeCommands;
			Sw12_state : in singleSwitchStates;
			Sw12_lock : in objectLock;
			Sw12_command : out routeCommands;
			Sw13_state : in singleSwitchStates;
			Sw13_lock : in objectLock;
			Sw13_command : out routeCommands;
			S122_state : in signalStates;
			S122_lock : in objectLock;
			S122_command : out routeCommands;
			T21_state : in signalStates;
			routeState : out std_logic
		);
	end component route_75;
	component route_76 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne41_state : in nodeStates;
			ne41_lock : in objectLock;
			ne41_command : out routeCommands;
			ne82_state : in nodeStates;
			ne82_lock : in objectLock;
			ne82_command : out routeCommands;
			ne32_state : in nodeStates;
			ne32_lock : in objectLock;
			ne32_command : out routeCommands;
			Sw04_state : in singleSwitchStates;
			Sw04_lock : in objectLock;
			Sw04_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			B130_state : in signalStates;
			B130_lock : in objectLock;
			B130_command : out routeCommands;
			C100_state : in signalStates;
			routeState : out std_logic
		);
	end component route_76;
	component route_77 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne41_state : in nodeStates;
			ne41_lock : in objectLock;
			ne41_command : out routeCommands;
			ne85_state : in nodeStates;
			ne85_lock : in objectLock;
			ne85_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			ne44_state : in nodeStates;
			ne44_lock : in objectLock;
			ne44_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			Sw41_state : in singleSwitchStates;
			Sw41_lock : in objectLock;
			Sw41_command : out routeCommands;
			B130_state : in signalStates;
			B130_lock : in objectLock;
			B130_command : out routeCommands;
			S105_state : in signalStates;
			routeState : out std_logic
		);
	end component route_77;
	component route_78 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne85_state : in nodeStates;
			ne85_lock : in objectLock;
			ne85_command : out routeCommands;
			ne41_state : in nodeStates;
			ne41_lock : in objectLock;
			ne41_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			S131_state : in signalStates;
			S131_lock : in objectLock;
			S131_command : out routeCommands;
			P58_state : in signalStates;
			routeState : out std_logic
		);
	end component route_78;
	component route_79 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne85_state : in nodeStates;
			ne85_lock : in objectLock;
			ne85_command : out routeCommands;
			ne84_state : in nodeStates;
			ne84_lock : in objectLock;
			ne84_command : out routeCommands;
			Sw05_state : in doubleSwitchStates;
			Sw05_lock : in objectLock;
			Sw05_command : out routeCommands;
			S131_state : in signalStates;
			S131_lock : in objectLock;
			S131_command : out routeCommands;
			T13_state : in signalStates;
			routeState : out std_logic
		);
	end component route_79;
	component route_80 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne77_state : in nodeStates;
			ne77_lock : in objectLock;
			ne77_command : out routeCommands;
			ne52_state : in nodeStates;
			ne52_lock : in objectLock;
			ne52_command : out routeCommands;
			Sw03_state : in scissorCrossingStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			B133_state : in signalStates;
			B133_lock : in objectLock;
			B133_command : out routeCommands;
			S86_state : in signalStates;
			routeState : out std_logic
		);
	end component route_80;
	component route_81 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne94_state : in nodeStates;
			ne94_lock : in objectLock;
			ne94_command : out routeCommands;
			ne77_state : in nodeStates;
			ne77_lock : in objectLock;
			ne77_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			S135_state : in signalStates;
			S135_lock : in objectLock;
			S135_command : out routeCommands;
			B133_state : in signalStates;
			routeState : out std_logic
		);
	end component route_81;
	component route_82 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne94_state : in nodeStates;
			ne94_lock : in objectLock;
			ne94_command : out routeCommands;
			ne21_state : in nodeStates;
			ne21_lock : in objectLock;
			ne21_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			S135_state : in signalStates;
			S135_lock : in objectLock;
			S135_command : out routeCommands;
			P72_state : in signalStates;
			routeState : out std_logic
		);
	end component route_82;
	component route_83 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			ne101_state : in nodeStates;
			ne101_lock : in objectLock;
			ne101_command : out routeCommands;
			ne44_state : in nodeStates;
			ne44_lock : in objectLock;
			ne44_command : out routeCommands;
			Sw41_state : in singleSwitchStates;
			Sw41_lock : in objectLock;
			Sw41_command : out routeCommands;
			C138_state : in signalStates;
			C138_lock : in objectLock;
			C138_command : out routeCommands;
			S105_state : in signalStates;
			routeState : out std_logic
		);
	end component route_83;
	component route_84 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			ne110_state : in nodeStates;
			ne110_lock : in objectLock;
			ne110_command : out routeCommands;
			Sw41_state : in singleSwitchStates;
			Sw41_lock : in objectLock;
			Sw41_command : out routeCommands;
			S139_state : in signalStates;
			S139_lock : in objectLock;
			S139_command : out routeCommands;
			S102_state : in signalStates;
			routeState : out std_logic
		);
	end component route_84;
	component route_85 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne100_state : in nodeStates;
			ne100_lock : in objectLock;
			ne100_command : out routeCommands;
			ne85_state : in nodeStates;
			ne85_lock : in objectLock;
			ne85_command : out routeCommands;
			Sw41_state : in singleSwitchStates;
			Sw41_lock : in objectLock;
			Sw41_command : out routeCommands;
			S139_state : in signalStates;
			S139_lock : in objectLock;
			S139_command : out routeCommands;
			S131_state : in signalStates;
			routeState : out std_logic
		);
	end component route_85;
	component route_86 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne104_state : in nodeStates;
			ne104_lock : in objectLock;
			ne104_command : out routeCommands;
			ne70_state : in nodeStates;
			ne70_lock : in objectLock;
			ne70_command : out routeCommands;
			B143_state : in signalStates;
			B143_lock : in objectLock;
			B143_command : out routeCommands;
			L32_state : in signalStates;
			routeState : out std_logic
		);
	end component route_86;
	component route_87 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne21_state : in nodeStates;
			ne21_lock : in objectLock;
			ne21_command : out routeCommands;
			ne104_state : in nodeStates;
			ne104_lock : in objectLock;
			ne104_command : out routeCommands;
			Sw03_state : in scissorCrossingStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			S144_state : in signalStates;
			S144_lock : in objectLock;
			S144_command : out routeCommands;
			B143_state : in signalStates;
			routeState : out std_logic
		);
	end component route_87;
	component route_88 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne77_state : in nodeStates;
			ne77_lock : in objectLock;
			ne77_command : out routeCommands;
			ne79_state : in nodeStates;
			ne79_lock : in objectLock;
			ne79_command : out routeCommands;
			ne78_state : in nodeStates;
			ne78_lock : in objectLock;
			ne78_command : out routeCommands;
			Sw06_state : in singleSwitchStates;
			Sw06_lock : in objectLock;
			Sw06_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			B145_state : in signalStates;
			B145_lock : in objectLock;
			B145_command : out routeCommands;
			L33_state : in signalStates;
			routeState : out std_logic
		);
	end component route_88;
	component route_89 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne77_state : in nodeStates;
			ne77_lock : in objectLock;
			ne77_command : out routeCommands;
			ne94_state : in nodeStates;
			ne94_lock : in objectLock;
			ne94_command : out routeCommands;
			ne97_state : in nodeStates;
			ne97_lock : in objectLock;
			ne97_command : out routeCommands;
			ne99_state : in nodeStates;
			ne99_lock : in objectLock;
			ne99_command : out routeCommands;
			Sw07_state : in doubleSwitchStates;
			Sw07_lock : in objectLock;
			Sw07_command : out routeCommands;
			B145_state : in signalStates;
			B145_lock : in objectLock;
			B145_command : out routeCommands;
			P69_state : in signalStates;
			routeState : out std_logic
		);
	end component route_89;
	component route_90 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			routeRequest : in std_logic;
			ne52_state : in nodeStates;
			ne52_lock : in objectLock;
			ne52_command : out routeCommands;
			ne77_state : in nodeStates;
			ne77_lock : in objectLock;
			ne77_command : out routeCommands;
			Sw03_state : in scissorCrossingStates;
			Sw03_lock : in objectLock;
			Sw03_command : out routeCommands;
			S146_state : in signalStates;
			S146_lock : in objectLock;
			S146_command : out routeCommands;
			B145_state : in signalStates;
			routeState : out std_logic
		);
	end component route_90;
	signal state_Lc01 : levelCrossingStates;
	signal Lc01_locking : objectLock;
	signal state_68W02 , state_69W03 , state_69W04 , state_Sw06 , state_70W01 , state_70W02 , state_Sw08 , state_Sw09 , state_Sw12 , state_Sw04 , state_71W01 , state_71W02 , state_Sw11 , state_Sw13 , state_Sw41 : singleSwitchStates;
	signal s68W02_locking , s69W03_locking , s69W04_locking , Sw06_locking , s70W01_locking , s70W02_locking , Sw08_locking , Sw09_locking , Sw12_locking , Sw04_locking , s71W01_locking , s71W02_locking , Sw11_locking , Sw13_locking , Sw41_locking : objectLock;
	signal state_Sw03 : scissorCrossingStates;
	signal Sw03_locking : objectLock;
	signal state_Sw05 , state_Sw07 : doubleSwitchStates;
	signal Sw05_locking , Sw07_locking : objectLock;
	signal state_T01 , state_T02 , state_C78 , state_T03 , state_L25 , state_T05 , state_T06 , state_J43 , state_J46 , state_S80 , state_T07 , state_T08 , state_C82 , state_C109 , state_P60 , state_B89 , state_P63 , state_B92 , state_L27 , state_S93 , state_B96 , state_B101 , state_S97 , state_S122 , state_C100 , state_S115 , state_P58 , state_B130 , state_L28 , state_S105 , state_T11 , state_T12 , state_L29 , state_S83 , state_S90 , state_L30 , state_P64 , state_P65 , state_L32 , state_L33 , state_S110 , state_C95 , state_C114 , state_T13 , state_T14 , state_T15 , state_S119 , state_T17 , state_C118 , state_T19 , state_T20 , state_T21 , state_T22 , state_L34 , state_S135 , state_L35 , state_X50 , state_X51 , state_P70 , state_P71 , state_L37 , state_L38 , state_P68 , state_P69 , state_S139 , state_L40 , state_C104 , state_L41 , state_T23 , state_T24 , state_L42 , state_S131 , state_B133 , state_B145 , state_B143 , state_S86 , state_S146 , state_P72 , state_P73 , state_S144 , state_S102 , state_C138 : signalStates;
	signal T01_locking , T02_locking , C78_locking , T03_locking , L25_locking , T05_locking , T06_locking , J43_locking , J46_locking , S80_locking , T07_locking , T08_locking , C82_locking , C109_locking , P60_locking , B89_locking , P63_locking , B92_locking , L27_locking , S93_locking , B96_locking , B101_locking , S97_locking , S122_locking , C100_locking , S115_locking , P58_locking , B130_locking , L28_locking , S105_locking , T11_locking , T12_locking , L29_locking , S83_locking , S90_locking , L30_locking , P64_locking , P65_locking , L32_locking , L33_locking , S110_locking , C95_locking , C114_locking , T13_locking , T14_locking , T15_locking , S119_locking , T17_locking , C118_locking , T19_locking , T20_locking , T21_locking , T22_locking , L34_locking , S135_locking , L35_locking , X50_locking , X51_locking , P70_locking , P71_locking , L37_locking , L38_locking , P68_locking , P69_locking , S139_locking , L40_locking , C104_locking , L41_locking , T23_locking , T24_locking , L42_locking , S131_locking , B133_locking , B145_locking , B143_locking , S86_locking , S146_locking , P72_locking , P73_locking , S144_locking , S102_locking , C138_locking : objectLock;
	signal state_ne1 , state_ne4 , state_ne7 , state_ne9 , state_ne11 , state_ne14 , state_ne17 , state_ne23 , state_ne24 , state_ne26 , state_ne29 , state_ne30 , state_ne32 , state_ne41 , state_ne43 , state_ne44 , state_ne47 , state_ne48 , state_ne59 , state_ne64 , state_ne65 , state_ne67 , state_ne70 , state_ne78 , state_ne79 , state_ne82 , state_ne83 , state_ne84 , state_ne86 , state_ne87 , state_ne88 , state_ne89 , state_ne90 , state_ne91 , state_ne93 , state_ne94 , state_ne95 , state_ne96 , state_ne97 , state_ne98 , state_ne99 , state_ne100 , state_ne101 , state_ne102 , state_ne103 , state_ne105 , state_ne106 , state_ne85 , state_ne77 , state_ne104 , state_ne52 , state_ne21 , state_ne110 : nodeStates;
	signal ne1_locking , ne4_locking , ne7_locking , ne9_locking , ne11_locking , ne14_locking , ne17_locking , ne23_locking , ne24_locking , ne26_locking , ne29_locking , ne30_locking , ne32_locking , ne41_locking , ne43_locking , ne44_locking , ne47_locking , ne48_locking , ne59_locking , ne64_locking , ne65_locking , ne67_locking , ne70_locking , ne78_locking , ne79_locking , ne82_locking , ne83_locking , ne84_locking , ne86_locking , ne87_locking , ne88_locking , ne89_locking , ne90_locking , ne91_locking , ne93_locking , ne94_locking , ne95_locking , ne96_locking , ne97_locking , ne98_locking , ne99_locking , ne100_locking , ne101_locking , ne102_locking , ne103_locking , ne105_locking , ne106_locking , ne85_locking , ne77_locking , ne104_locking , ne52_locking , ne21_locking , ne110_locking : objectLock;
	signal cmd_R1_ne1 , cmd_R2_ne7 , cmd_R3_ne14 , cmd_R3_ne52 , cmd_R4_ne47 , cmd_R4_ne48 , cmd_R5_ne84 , cmd_R5_ne82 , cmd_R5_ne32 , cmd_R6_ne84 , cmd_R6_ne85 , cmd_R6_ne100 , cmd_R6_ne101 , cmd_R6_ne44 , cmd_R7_ne89 , cmd_R7_ne30 , cmd_R8_ne90 , cmd_R8_ne91 , cmd_R8_ne30 , cmd_R9_ne105 , cmd_R9_ne98 , cmd_R9_ne96 , cmd_R10_ne4 , cmd_R10_ne106 , cmd_R11_ne26 , cmd_R11_ne65 , cmd_R12_ne44 , cmd_R12_ne101 , cmd_R13_ne65 , cmd_R13_ne102 , cmd_R14_ne70 , cmd_R14_ne104 , cmd_R14_ne21 , cmd_R15_ne78 , cmd_R15_ne93 , cmd_R16_ne93 , cmd_R16_ne96 , cmd_R17_ne95 , cmd_R18_ne97 , cmd_R18_ne94 , cmd_R19_ne98 , cmd_R19_ne105 , cmd_R20_ne101 , cmd_R20_ne100 , cmd_R21_ne103 , cmd_R21_ne64 , cmd_R22_ne106 , cmd_R22_ne99 , cmd_R23_ne7 , cmd_R23_ne9 , cmd_R24_ne9 , cmd_R24_ne95 , cmd_R25_ne95 , cmd_R25_ne59 , cmd_R26_ne95 , cmd_R26_ne9 , cmd_R27_ne23 , cmd_R27_ne26 , cmd_R28_ne24 , cmd_R28_ne64 , cmd_R28_ne103 , cmd_R28_ne67 , cmd_R29_ne67 , cmd_R29_ne70 , cmd_R30_ne67 , cmd_R30_ne103 , cmd_R31_ne99 , cmd_R31_ne97 , cmd_R32_ne99 , cmd_R32_ne106 , cmd_R32_ne4 , cmd_R33_ne96 , cmd_R33_ne93 , cmd_R33_ne78 , cmd_R34_ne96 , cmd_R34_ne98 , cmd_R35_ne21 , cmd_R36_ne21 , cmd_R36_ne79 , cmd_R36_ne78 , cmd_R37_ne21 , cmd_R37_ne94 , cmd_R37_ne97 , cmd_R37_ne99 , cmd_R38_ne1 , cmd_R38_ne9 , cmd_R39_ne9 , cmd_R39_ne1 , cmd_R40_ne9 , cmd_R40_ne7 , cmd_R41_ne17 , cmd_R41_ne59 , cmd_R41_ne95 , cmd_R42_ne59 , cmd_R42_ne11 , cmd_R42_ne52 , cmd_R43_ne59 , cmd_R43_ne17 , cmd_R44_ne52 , cmd_R44_ne11 , cmd_R44_ne59 , cmd_R44_ne95 , cmd_R45_ne52 , cmd_R45_ne14 , cmd_R46_ne23 , cmd_R46_ne64 , cmd_R46_ne103 , cmd_R46_ne67 , cmd_R47_ne64 , cmd_R47_ne23 , cmd_R48_ne64 , cmd_R48_ne24 , cmd_R49_ne24 , cmd_R49_ne26 , cmd_R50_ne26 , cmd_R50_ne23 , cmd_R51_ne26 , cmd_R51_ne24 , cmd_R52_ne83 , cmd_R52_ne30 , cmd_R53_ne29 , cmd_R53_ne30 , cmd_R54_ne30 , cmd_R54_ne29 , cmd_R54_ne110 , cmd_R55_ne30 , cmd_R55_ne83 , cmd_R56_ne32 , cmd_R56_ne110 , cmd_R57_ne29 , cmd_R58_ne110 , cmd_R58_ne32 , cmd_R59_ne110 , cmd_R59_ne29 , cmd_R60_ne102 , cmd_R60_ne44 , cmd_R61_ne44 , cmd_R61_ne43 , cmd_R61_ne48 , cmd_R62_ne44 , cmd_R62_ne102 , cmd_R62_ne65 , cmd_R62_ne26 , cmd_R63_ne17 , cmd_R63_ne78 , cmd_R64_ne78 , cmd_R64_ne17 , cmd_R65_ne78 , cmd_R65_ne79 , cmd_R65_ne77 , cmd_R66_ne78 , cmd_R66_ne79 , cmd_R66_ne21 , cmd_R67_ne83 , cmd_R67_ne32 , cmd_R68_ne32 , cmd_R68_ne83 , cmd_R69_ne32 , cmd_R69_ne82 , cmd_R69_ne41 , cmd_R70_ne32 , cmd_R70_ne82 , cmd_R70_ne84 , cmd_R71_ne88 , cmd_R71_ne86 , cmd_R72_ne86 , cmd_R72_ne88 , cmd_R73_ne86 , cmd_R73_ne87 , cmd_R73_ne91 , cmd_R73_ne30 , cmd_R74_ne30 , cmd_R74_ne89 , cmd_R75_ne30 , cmd_R75_ne91 , cmd_R75_ne87 , cmd_R75_ne86 , cmd_R76_ne30 , cmd_R76_ne91 , cmd_R76_ne90 , cmd_R77_ne41 , cmd_R77_ne82 , cmd_R77_ne32 , cmd_R78_ne41 , cmd_R78_ne85 , cmd_R78_ne100 , cmd_R78_ne101 , cmd_R78_ne44 , cmd_R79_ne85 , cmd_R79_ne41 , cmd_R80_ne85 , cmd_R80_ne84 , cmd_R81_ne77 , cmd_R81_ne52 , cmd_R82_ne94 , cmd_R82_ne77 , cmd_R83_ne94 , cmd_R83_ne21 , cmd_R84_ne110 , cmd_R84_ne100 , cmd_R84_ne101 , cmd_R84_ne44 , cmd_R85_ne100 , cmd_R85_ne110 , cmd_R86_ne100 , cmd_R86_ne85 , cmd_R87_ne104 , cmd_R87_ne70 , cmd_R88_ne21 , cmd_R88_ne104 , cmd_R89_ne77 , cmd_R89_ne79 , cmd_R89_ne78 , cmd_R90_ne77 , cmd_R90_ne94 , cmd_R90_ne97 , cmd_R90_ne99 , cmd_R91_ne52 , cmd_R91_ne77 : routeCommands;
	signal cmd_R25_Lc01 , cmd_R26_Lc01 : routeCommands;
	signal cmd_R3_69W04 , cmd_R4_71W02 , cmd_R5_Sw04 , cmd_R5_Sw05 , cmd_R6_Sw05 , cmd_R6_Sw41 , cmd_R7_Sw12 , cmd_R8_Sw12 , cmd_R8_Sw13 , cmd_R23_68W02 , cmd_R27_70W02 , cmd_R36_Sw06 , cmd_R36_Sw07 , cmd_R37_Sw07 , cmd_R38_68W02 , cmd_R39_68W02 , cmd_R40_68W02 , cmd_R41_69W03 , cmd_R42_69W03 , cmd_R42_69W04 , cmd_R43_69W03 , cmd_R44_69W03 , cmd_R44_69W04 , cmd_R45_69W04 , cmd_R47_70W01 , cmd_R48_70W01 , cmd_R49_70W02 , cmd_R50_70W02 , cmd_R51_70W02 , cmd_R52_Sw08 , cmd_R53_Sw08 , cmd_R54_Sw08 , cmd_R54_Sw09 , cmd_R55_Sw08 , cmd_R56_Sw09 , cmd_R58_Sw09 , cmd_R59_Sw09 , cmd_R60_71W01 , cmd_R61_71W01 , cmd_R61_71W02 , cmd_R62_71W01 , cmd_R63_Sw06 , cmd_R64_Sw06 , cmd_R65_Sw06 , cmd_R65_Sw07 , cmd_R66_Sw06 , cmd_R66_Sw07 , cmd_R67_Sw04 , cmd_R68_Sw04 , cmd_R69_Sw04 , cmd_R69_Sw05 , cmd_R70_Sw04 , cmd_R70_Sw05 , cmd_R71_Sw11 , cmd_R72_Sw11 , cmd_R73_Sw11 , cmd_R73_Sw12 , cmd_R73_Sw13 , cmd_R74_Sw12 , cmd_R75_Sw11 , cmd_R75_Sw12 , cmd_R75_Sw13 , cmd_R76_Sw12 , cmd_R76_Sw13 , cmd_R77_Sw04 , cmd_R77_Sw05 , cmd_R78_Sw05 , cmd_R78_Sw41 , cmd_R79_Sw05 , cmd_R80_Sw05 , cmd_R82_Sw07 , cmd_R83_Sw07 , cmd_R84_Sw41 , cmd_R85_Sw41 , cmd_R86_Sw41 , cmd_R89_Sw06 , cmd_R89_Sw07 , cmd_R90_Sw07 : routeCommands;
	signal cmd_R14_Sw03 , cmd_R81_Sw03 , cmd_R88_Sw03 , cmd_R91_Sw03 : routeCommands;
	signal cmd_R1_T02 , cmd_R2_T06 , cmd_R3_T08 , cmd_R4_T12 , cmd_R5_T14 , cmd_R6_T14 , cmd_R7_T20 , cmd_R8_T22 , cmd_R9_T24 , cmd_R10_L25 , cmd_R11_L27 , cmd_R12_L28 , cmd_R13_L30 , cmd_R14_L32 , cmd_R15_L33 , cmd_R16_L34 , cmd_R17_L35 , cmd_R18_L37 , cmd_R19_L38 , cmd_R20_L40 , cmd_R21_L41 , cmd_R22_L42 , cmd_R23_J43 , cmd_R24_J46 , cmd_R25_X50 , cmd_R26_X51 , cmd_R27_P60 , cmd_R28_P63 , cmd_R29_P64 , cmd_R30_P65 , cmd_R31_P68 , cmd_R32_P69 , cmd_R33_P70 , cmd_R34_P71 , cmd_R35_P72 , cmd_R36_P73 , cmd_R37_P73 , cmd_R38_C78 , cmd_R39_S80 , cmd_R40_S80 , cmd_R41_C82 , cmd_R42_S83 , cmd_R43_S83 , cmd_R44_S86 , cmd_R45_S86 , cmd_R46_B89 , cmd_R47_S90 , cmd_R48_S90 , cmd_R49_B92 , cmd_R50_S93 , cmd_R51_S93 , cmd_R52_C95 , cmd_R53_B96 , cmd_R54_S97 , cmd_R55_S97 , cmd_R56_C100 , cmd_R57_B101 , cmd_R58_S102 , cmd_R59_S102 , cmd_R60_C104 , cmd_R61_S105 , cmd_R62_S105 , cmd_R63_C109 , cmd_R64_S110 , cmd_R65_S110 , cmd_R66_S110 , cmd_R67_C114 , cmd_R68_S115 , cmd_R69_S115 , cmd_R70_S115 , cmd_R71_C118 , cmd_R72_S119 , cmd_R73_S119 , cmd_R74_S122 , cmd_R75_S122 , cmd_R76_S122 , cmd_R77_B130 , cmd_R78_B130 , cmd_R79_S131 , cmd_R80_S131 , cmd_R81_B133 , cmd_R82_S135 , cmd_R83_S135 , cmd_R84_C138 , cmd_R85_S139 , cmd_R86_S139 , cmd_R87_B143 , cmd_R88_S144 , cmd_R89_B145 , cmd_R90_B145 , cmd_R91_S146 : routeCommands;
begin
	levelCrossing_Lc01 : levelCrossing_0 port map(clock => clock, reset => reset, R25_command => cmd_R25_Lc01, R26_command => cmd_R26_Lc01, ocupation_ne95 => ocupation(36), ocupation_ne9 => ocupation(3), ocupation_ne59 => ocupation(18), indication => levelCrossings_i, command  => levelCrossings_o, lock_Lc01 => Lc01_locking, correspondence_Lc01 => state_Lc01);
	singleSwitch_68W02 : singleSwitch_0 port map(clock => clock, reset => reset, R23_command => cmd_R23_68W02, R38_command => cmd_R38_68W02, R39_command => cmd_R39_68W02, R40_command => cmd_R40_68W02, indication => singleSwitches_i(0), command => singleSwitches_o(0), lock_68W02 => s68W02_locking, correspondence_68W02 => state_68W02);
	singleSwitch_69W03 : singleSwitch_1 port map(clock => clock, reset => reset, R41_command => cmd_R41_69W03, R42_command => cmd_R42_69W03, R43_command => cmd_R43_69W03, R44_command => cmd_R44_69W03, indication => singleSwitches_i(1), command => singleSwitches_o(1), lock_69W03 => s69W03_locking, correspondence_69W03 => state_69W03);
	singleSwitch_69W04 : singleSwitch_2 port map(clock => clock, reset => reset, R3_command => cmd_R3_69W04, R42_command => cmd_R42_69W04, R44_command => cmd_R44_69W04, R45_command => cmd_R45_69W04, indication => singleSwitches_i(2), command => singleSwitches_o(2), lock_69W04 => s69W04_locking, correspondence_69W04 => state_69W04);
	singleSwitch_Sw06 : singleSwitch_3 port map(clock => clock, reset => reset, R36_command => cmd_R36_Sw06, R63_command => cmd_R63_Sw06, R64_command => cmd_R64_Sw06, R65_command => cmd_R65_Sw06, R66_command => cmd_R66_Sw06, R89_command => cmd_R89_Sw06, indication => singleSwitches_i(3), command => singleSwitches_o(3), lock_Sw06 => Sw06_locking, correspondence_Sw06 => state_Sw06);
	singleSwitch_70W01 : singleSwitch_4 port map(clock => clock, reset => reset, R47_command => cmd_R47_70W01, R48_command => cmd_R48_70W01, indication => singleSwitches_i(4), command => singleSwitches_o(4), lock_70W01 => s70W01_locking, correspondence_70W01 => state_70W01);
	singleSwitch_70W02 : singleSwitch_5 port map(clock => clock, reset => reset, R27_command => cmd_R27_70W02, R49_command => cmd_R49_70W02, R50_command => cmd_R50_70W02, R51_command => cmd_R51_70W02, indication => singleSwitches_i(5), command => singleSwitches_o(5), lock_70W02 => s70W02_locking, correspondence_70W02 => state_70W02);
	singleSwitch_Sw08 : singleSwitch_6 port map(clock => clock, reset => reset, R52_command => cmd_R52_Sw08, R53_command => cmd_R53_Sw08, R54_command => cmd_R54_Sw08, R55_command => cmd_R55_Sw08, indication => singleSwitches_i(6), command => singleSwitches_o(6), lock_Sw08 => Sw08_locking, correspondence_Sw08 => state_Sw08);
	singleSwitch_Sw09 : singleSwitch_7 port map(clock => clock, reset => reset, R54_command => cmd_R54_Sw09, R56_command => cmd_R56_Sw09, R58_command => cmd_R58_Sw09, R59_command => cmd_R59_Sw09, indication => singleSwitches_i(7), command => singleSwitches_o(7), lock_Sw09 => Sw09_locking, correspondence_Sw09 => state_Sw09);
	singleSwitch_Sw12 : singleSwitch_8 port map(clock => clock, reset => reset, R7_command => cmd_R7_Sw12, R8_command => cmd_R8_Sw12, R73_command => cmd_R73_Sw12, R74_command => cmd_R74_Sw12, R75_command => cmd_R75_Sw12, R76_command => cmd_R76_Sw12, indication => singleSwitches_i(8), command => singleSwitches_o(8), lock_Sw12 => Sw12_locking, correspondence_Sw12 => state_Sw12);
	singleSwitch_Sw04 : singleSwitch_9 port map(clock => clock, reset => reset, R5_command => cmd_R5_Sw04, R67_command => cmd_R67_Sw04, R68_command => cmd_R68_Sw04, R69_command => cmd_R69_Sw04, R70_command => cmd_R70_Sw04, R77_command => cmd_R77_Sw04, indication => singleSwitches_i(9), command => singleSwitches_o(9), lock_Sw04 => Sw04_locking, correspondence_Sw04 => state_Sw04);
	singleSwitch_71W01 : singleSwitch_10 port map(clock => clock, reset => reset, R60_command => cmd_R60_71W01, R61_command => cmd_R61_71W01, R62_command => cmd_R62_71W01, indication => singleSwitches_i(10), command => singleSwitches_o(10), lock_71W01 => s71W01_locking, correspondence_71W01 => state_71W01);
	singleSwitch_71W02 : singleSwitch_11 port map(clock => clock, reset => reset, R4_command => cmd_R4_71W02, R61_command => cmd_R61_71W02, indication => singleSwitches_i(11), command => singleSwitches_o(11), lock_71W02 => s71W02_locking, correspondence_71W02 => state_71W02);
	singleSwitch_Sw11 : singleSwitch_12 port map(clock => clock, reset => reset, R71_command => cmd_R71_Sw11, R72_command => cmd_R72_Sw11, R73_command => cmd_R73_Sw11, R75_command => cmd_R75_Sw11, indication => singleSwitches_i(12), command => singleSwitches_o(12), lock_Sw11 => Sw11_locking, correspondence_Sw11 => state_Sw11);
	singleSwitch_Sw13 : singleSwitch_13 port map(clock => clock, reset => reset, R8_command => cmd_R8_Sw13, R73_command => cmd_R73_Sw13, R75_command => cmd_R75_Sw13, R76_command => cmd_R76_Sw13, indication => singleSwitches_i(13), command => singleSwitches_o(13), lock_Sw13 => Sw13_locking, correspondence_Sw13 => state_Sw13);
	singleSwitch_Sw41 : singleSwitch_14 port map(clock => clock, reset => reset, R6_command => cmd_R6_Sw41, R78_command => cmd_R78_Sw41, R84_command => cmd_R84_Sw41, R85_command => cmd_R85_Sw41, R86_command => cmd_R86_Sw41, indication => singleSwitches_i(14), command => singleSwitches_o(14), lock_Sw41 => Sw41_locking, correspondence_Sw41 => state_Sw41);
	scissorCrossing_Sw03 : scissorCrossing_0 port map(clock => clock, reset => reset, R14_command => cmd_R14_Sw03, R81_command => cmd_R81_Sw03, R88_command => cmd_R88_Sw03, R91_command => cmd_R91_Sw03, indication => scissorCrossings_i, command => scissorCrossings_o, lock_Sw03 => Sw03_locking, correspondence_Sw03 => state_Sw03);
	doubleSwitch_Sw05 : doubleSwitch_0 port map(clock => clock, reset => reset, R5_command => cmd_R5_Sw05, R6_command => cmd_R6_Sw05, R69_command => cmd_R69_Sw05, R70_command => cmd_R70_Sw05, R77_command => cmd_R77_Sw05, R78_command => cmd_R78_Sw05, R79_command => cmd_R79_Sw05, R80_command => cmd_R80_Sw05, indication.msb => doubleSwitches_i.msb(0), indication.lsb => doubleSwitches_i.lsb(0), command.msb => doubleSwitches_o.msb(0), command.lsb => doubleSwitches_o.lsb(0),lock_Sw05 => Sw05_locking, correspondence_Sw05 => state_Sw05);
	doubleSwitch_Sw07 : doubleSwitch_1 port map(clock => clock, reset => reset, R36_command => cmd_R36_Sw07, R37_command => cmd_R37_Sw07, R65_command => cmd_R65_Sw07, R66_command => cmd_R66_Sw07, R82_command => cmd_R82_Sw07, R83_command => cmd_R83_Sw07, R89_command => cmd_R89_Sw07, R90_command => cmd_R90_Sw07, indication.msb => doubleSwitches_i.msb(1), indication.lsb => doubleSwitches_i.lsb(1), command.msb => doubleSwitches_o.msb(1), command.lsb => doubleSwitches_o.lsb(1),lock_Sw07 => Sw07_locking, correspondence_Sw07 => state_Sw07);
	railwaySignal_T01 : railwaySignal_0 port map(clock => clock, reset => reset, ocupation_ne1 => ocupation(0), indication.msb => signals_i.msb(0), indication.lsb => signals_i.lsb(0), command.msb => signals_o.msb(0), command.lsb => signals_o.lsb(0), lock_T01 => T01_locking, correspondence_T01 => state_T01);
	railwaySignal_T02 : railwaySignal_1 port map(clock => clock, reset => reset, R1_command => cmd_R1_T02, ocupation_ne1 => ocupation(0), ocupation_ne9 => ocupation(3), correspondence_C78 => state_C78, correspondence_J46 => state_J46, s68W02_state => state_68W02, indication.msb => signals_i.msb(1), indication.lsb => signals_i.lsb(1), command.msb => signals_o.msb(1), command.lsb => signals_o.lsb(1), lock_T02 => T02_locking, correspondence_T02 => state_T02);
	railwaySignal_C78 : railwaySignal_2 port map(clock => clock, reset => reset, R38_command => cmd_R38_C78, ocupation_ne1 => ocupation(0), ocupation_ne9 => ocupation(3), ocupation_ne95 => ocupation(36), correspondence_J46 => state_J46, correspondence_L35 => state_L35, s68W02_state => state_68W02, indication.msb => signals_i.msb(2), indication.lsb => signals_i.lsb(2), command.msb => signals_o.msb(2), command.lsb => signals_o.lsb(2), lock_C78 => C78_locking, correspondence_C78 => state_C78);
	railwaySignal_T03 : railwaySignal_3 port map(clock => clock, reset => reset, ocupation_ne4 => ocupation(1), indication.msb => signals_i.msb(3), indication.lsb => signals_i.lsb(3), command.msb => signals_o.msb(3), command.lsb => signals_o.lsb(3), lock_T03 => T03_locking, correspondence_T03 => state_T03);
	railwaySignal_L25 : railwaySignal_4 port map(clock => clock, reset => reset, R10_command => cmd_R10_L25, ocupation_ne4 => ocupation(1), ocupation_ne106 => ocupation(46), ocupation_ne99 => ocupation(40), correspondence_L42 => state_L42, correspondence_P68 => state_P68, indication.msb => signals_i.msb(4), indication.lsb => signals_i.lsb(4), command.msb => signals_o.msb(4), command.lsb => signals_o.lsb(4), lock_L25 => L25_locking, correspondence_L25 => state_L25);
	railwaySignal_T05 : railwaySignal_5 port map(clock => clock, reset => reset, ocupation_ne7 => ocupation(2), indication.msb => signals_i.msb(5), indication.lsb => signals_i.lsb(5), command.msb => signals_o.msb(5), command.lsb => signals_o.lsb(5), lock_T05 => T05_locking, correspondence_T05 => state_T05);
	railwaySignal_T06 : railwaySignal_6 port map(clock => clock, reset => reset, R2_command => cmd_R2_T06, ocupation_ne7 => ocupation(2), ocupation_ne9 => ocupation(3), correspondence_J43 => state_J43, correspondence_J46 => state_J46, s68W02_state => state_68W02, indication.msb => signals_i.msb(6), indication.lsb => signals_i.lsb(6), command.msb => signals_o.msb(6), command.lsb => signals_o.lsb(6), lock_T06 => T06_locking, correspondence_T06 => state_T06);
	railwaySignal_J43 : railwaySignal_7 port map(clock => clock, reset => reset, R23_command => cmd_R23_J43, ocupation_ne7 => ocupation(2), ocupation_ne9 => ocupation(3), ocupation_ne95 => ocupation(36), correspondence_J46 => state_J46, correspondence_L35 => state_L35, s68W02_state => state_68W02, indication.msb => signals_i.msb(7), indication.lsb => signals_i.lsb(7), command.msb => signals_o.msb(7), command.lsb => signals_o.lsb(7), lock_J43 => J43_locking, correspondence_J43 => state_J43);
	railwaySignal_J46 : railwaySignal_8 port map(clock => clock, reset => reset, R24_command => cmd_R24_J46, ocupation_ne9 => ocupation(3), ocupation_ne95 => ocupation(36), correspondence_L35 => state_L35, correspondence_X50 => state_X50, indication.msb => signals_i.msb(8), indication.lsb => signals_i.lsb(8), command.msb => signals_o.msb(8), command.lsb => signals_o.lsb(8), lock_J46 => J46_locking, correspondence_J46 => state_J46);
	railwaySignal_S80 : railwaySignal_9 port map(clock => clock, reset => reset, R39_command => cmd_R39_S80, R40_command => cmd_R40_S80, ocupation_ne9 => ocupation(3), ocupation_ne1 => ocupation(0), ocupation_ne7 => ocupation(2), correspondence_T01 => state_T01, correspondence_T05 => state_T05, s68W02_state => state_68W02, indication.msb => signals_i.msb(9), indication.lsb => signals_i.lsb(9), command.msb => signals_o.msb(9), command.lsb => signals_o.lsb(9), lock_S80 => S80_locking, correspondence_S80 => state_S80);
	railwaySignal_T07 : railwaySignal_10 port map(clock => clock, reset => reset, ocupation_ne14 => ocupation(5), indication.msb => signals_i.msb(10), indication.lsb => signals_i.lsb(10), command.msb => signals_o.msb(10), command.lsb => signals_o.lsb(10), lock_T07 => T07_locking, correspondence_T07 => state_T07);
	railwaySignal_T08 : railwaySignal_11 port map(clock => clock, reset => reset, R3_command => cmd_R3_T08, ocupation_ne14 => ocupation(5), ocupation_ne52 => ocupation(50), ocupation_ne77 => ocupation(48), correspondence_S146 => state_S146, correspondence_B145 => state_B145, s69W04_state => state_69W04, Sw03_state => state_Sw03, indication.msb => signals_i.msb(11), indication.lsb => signals_i.lsb(11), command.msb => signals_o.msb(11), command.lsb => signals_o.lsb(11), lock_T08 => T08_locking, correspondence_T08 => state_T08);
	railwaySignal_C82 : railwaySignal_12 port map(clock => clock, reset => reset, R41_command => cmd_R41_C82, ocupation_ne17 => ocupation(6), ocupation_ne59 => ocupation(18), ocupation_ne95 => ocupation(36), ocupation_ne9 => ocupation(3), correspondence_X51 => state_X51, correspondence_S80 => state_S80, s69W03_state => state_69W03, Lc01_state => state_Lc01, indication.msb => signals_i.msb(12), indication.lsb => signals_i.lsb(12), command.msb => signals_o.msb(12), command.lsb => signals_o.lsb(12), lock_C82 => C82_locking, correspondence_C82 => state_C82);
	railwaySignal_C109 : railwaySignal_13 port map(clock => clock, reset => reset, R63_command => cmd_R63_C109, ocupation_ne17 => ocupation(6), ocupation_ne78 => ocupation(23), ocupation_ne93 => ocupation(34), correspondence_L33 => state_L33, correspondence_L34 => state_L34, Sw06_state => state_Sw06, indication.msb => signals_i.msb(13), indication.lsb => signals_i.lsb(13), command.msb => signals_o.msb(13), command.lsb => signals_o.lsb(13), lock_C109 => C109_locking, correspondence_C109 => state_C109);
	railwaySignal_P60 : railwaySignal_14 port map(clock => clock, reset => reset, R27_command => cmd_R27_P60, ocupation_ne23 => ocupation(7), ocupation_ne26 => ocupation(9), ocupation_ne65 => ocupation(20), correspondence_L27 => state_L27, correspondence_L30 => state_L30, s70W02_state => state_70W02, indication.msb => signals_i.msb(14), indication.lsb => signals_i.lsb(14), command.msb => signals_o.msb(14), command.lsb => signals_o.lsb(14), lock_P60 => P60_locking, correspondence_P60 => state_P60);
	railwaySignal_B89 : railwaySignal_15 port map(clock => clock, reset => reset, R46_command => cmd_R46_B89, ocupation_ne23 => ocupation(7), ocupation_ne64 => ocupation(19), ocupation_ne103 => ocupation(44), ocupation_ne67 => ocupation(21), ocupation_ne70 => ocupation(22), correspondence_P64 => state_P64, correspondence_L32 => state_L32, indication.msb => signals_i.msb(15), indication.lsb => signals_i.lsb(15), command.msb => signals_o.msb(15), command.lsb => signals_o.lsb(15), lock_B89 => B89_locking, correspondence_B89 => state_B89);
	railwaySignal_P63 : railwaySignal_16 port map(clock => clock, reset => reset, R28_command => cmd_R28_P63, ocupation_ne24 => ocupation(8), ocupation_ne64 => ocupation(19), ocupation_ne103 => ocupation(44), ocupation_ne67 => ocupation(21), ocupation_ne70 => ocupation(22), correspondence_P64 => state_P64, correspondence_L32 => state_L32, indication.msb => signals_i.msb(16), indication.lsb => signals_i.lsb(16), command.msb => signals_o.msb(16), command.lsb => signals_o.lsb(16), lock_P63 => P63_locking, correspondence_P63 => state_P63);
	railwaySignal_B92 : railwaySignal_17 port map(clock => clock, reset => reset, R49_command => cmd_R49_B92, ocupation_ne24 => ocupation(8), ocupation_ne26 => ocupation(9), ocupation_ne65 => ocupation(20), correspondence_L27 => state_L27, correspondence_L30 => state_L30, s70W02_state => state_70W02, indication.msb => signals_i.msb(17), indication.lsb => signals_i.lsb(17), command.msb => signals_o.msb(17), command.lsb => signals_o.lsb(17), lock_B92 => B92_locking, correspondence_B92 => state_B92);
	railwaySignal_L27 : railwaySignal_18 port map(clock => clock, reset => reset, R11_command => cmd_R11_L27, ocupation_ne26 => ocupation(9), ocupation_ne65 => ocupation(20), ocupation_ne102 => ocupation(43), correspondence_L30 => state_L30, correspondence_C104 => state_C104, indication.msb => signals_i.msb(18), indication.lsb => signals_i.lsb(18), command.msb => signals_o.msb(18), command.lsb => signals_o.lsb(18), lock_L27 => L27_locking, correspondence_L27 => state_L27);
	railwaySignal_S93 : railwaySignal_19 port map(clock => clock, reset => reset, R50_command => cmd_R50_S93, R51_command => cmd_R51_S93, ocupation_ne26 => ocupation(9), ocupation_ne23 => ocupation(7), ocupation_ne24 => ocupation(8), ocupation_ne67 => ocupation(21), ocupation_ne103 => ocupation(44), ocupation_ne64 => ocupation(19), correspondence_B89 => state_B89, correspondence_P63 => state_P63, correspondence_P64 => state_P64, s70W02_state => state_70W02, indication.msb => signals_i.msb(19), indication.lsb => signals_i.lsb(19), command.msb => signals_o.msb(19), command.lsb => signals_o.lsb(19), lock_S93 => S93_locking, correspondence_S93 => state_S93);
	railwaySignal_B96 : railwaySignal_20 port map(clock => clock, reset => reset, R53_command => cmd_R53_B96, ocupation_ne29 => ocupation(10), ocupation_ne30 => ocupation(11), ocupation_ne90 => ocupation(32), ocupation_ne91 => ocupation(33), ocupation_ne86 => ocupation(28), ocupation_ne87 => ocupation(29), ocupation_ne89 => ocupation(31), correspondence_S122 => state_S122, correspondence_T19 => state_T19, correspondence_T15 => state_T15, correspondence_T21 => state_T21, Sw08_state => state_Sw08, Sw12_state => state_Sw12, Sw11_state => state_Sw11, Sw13_state => state_Sw13, indication.msb => signals_i.msb(20), indication.lsb => signals_i.lsb(20), command.msb => signals_o.msb(20), command.lsb => signals_o.lsb(20), lock_B96 => B96_locking, correspondence_B96 => state_B96);
	railwaySignal_B101 : railwaySignal_21 port map(clock => clock, reset => reset, R57_command => cmd_R57_B101, ocupation_ne29 => ocupation(10), ocupation_ne30 => ocupation(11), correspondence_B96 => state_B96, correspondence_S122 => state_S122, Sw08_state => state_Sw08, indication.msb => signals_i.msb(21), indication.lsb => signals_i.lsb(21), command.msb => signals_o.msb(21), command.lsb => signals_o.lsb(21), lock_B101 => B101_locking, correspondence_B101 => state_B101);
	railwaySignal_S97 : railwaySignal_22 port map(clock => clock, reset => reset, R54_command => cmd_R54_S97, R55_command => cmd_R55_S97, ocupation_ne30 => ocupation(11), ocupation_ne29 => ocupation(10), ocupation_ne110 => ocupation(52), ocupation_ne83 => ocupation(26), ocupation_ne101 => ocupation(42), ocupation_ne100 => ocupation(41), ocupation_ne44 => ocupation(15), ocupation_ne32 => ocupation(12), correspondence_C138 => state_C138, correspondence_C114 => state_C114, correspondence_S105 => state_S105, correspondence_C100 => state_C100, Sw08_state => state_Sw08, Sw09_state => state_Sw09, Sw41_state => state_Sw41, Sw04_state => state_Sw04, indication.msb => signals_i.msb(22), indication.lsb => signals_i.lsb(22), command.msb => signals_o.msb(22), command.lsb => signals_o.lsb(22), lock_S97 => S97_locking, correspondence_S97 => state_S97);
	railwaySignal_S122 : railwaySignal_23 port map(clock => clock, reset => reset, R74_command => cmd_R74_S122, R75_command => cmd_R75_S122, R76_command => cmd_R76_S122, ocupation_ne30 => ocupation(11), ocupation_ne89 => ocupation(31), ocupation_ne91 => ocupation(33), ocupation_ne87 => ocupation(29), ocupation_ne86 => ocupation(28), ocupation_ne90 => ocupation(32), correspondence_T19 => state_T19, correspondence_T15 => state_T15, correspondence_T21 => state_T21, Sw12_state => state_Sw12, Sw11_state => state_Sw11, Sw13_state => state_Sw13, indication.msb => signals_i.msb(23), indication.lsb => signals_i.lsb(23), command.msb => signals_o.msb(23), command.lsb => signals_o.lsb(23), lock_S122 => S122_locking, correspondence_S122 => state_S122);
	railwaySignal_C100 : railwaySignal_24 port map(clock => clock, reset => reset, R56_command => cmd_R56_C100, ocupation_ne32 => ocupation(12), ocupation_ne110 => ocupation(52), ocupation_ne101 => ocupation(42), ocupation_ne100 => ocupation(41), ocupation_ne44 => ocupation(15), correspondence_C138 => state_C138, correspondence_S105 => state_S105, Sw09_state => state_Sw09, Sw41_state => state_Sw41, indication.msb => signals_i.msb(24), indication.lsb => signals_i.lsb(24), command.msb => signals_o.msb(24), command.lsb => signals_o.lsb(24), lock_C100 => C100_locking, correspondence_C100 => state_C100);
	railwaySignal_S115 : railwaySignal_25 port map(clock => clock, reset => reset, R68_command => cmd_R68_S115, R69_command => cmd_R69_S115, R70_command => cmd_R70_S115, ocupation_ne32 => ocupation(12), ocupation_ne83 => ocupation(26), ocupation_ne82 => ocupation(25), ocupation_ne41 => ocupation(13), ocupation_ne84 => ocupation(27), ocupation_ne30 => ocupation(11), correspondence_C95 => state_C95, correspondence_P58 => state_P58, correspondence_T13 => state_T13, correspondence_S122 => state_S122, Sw04_state => state_Sw04, Sw08_state => state_Sw08, Sw05_state => state_Sw05, indication.msb => signals_i.msb(25), indication.lsb => signals_i.lsb(25), command.msb => signals_o.msb(25), command.lsb => signals_o.lsb(25), lock_S115 => S115_locking, correspondence_S115 => state_S115);
	railwaySignal_P58 : railwaySignal_26 port map(clock => clock, reset => reset, ocupation_ne41 => ocupation(13), indication.msb => signals_i.msb(26), indication.lsb => signals_i.lsb(26), command.msb => signals_o.msb(26), command.lsb => signals_o.lsb(26), lock_P58 => P58_locking, correspondence_P58 => state_P58);
	railwaySignal_B130 : railwaySignal_27 port map(clock => clock, reset => reset, R77_command => cmd_R77_B130, R78_command => cmd_R78_B130, ocupation_ne41 => ocupation(13), ocupation_ne82 => ocupation(25), ocupation_ne32 => ocupation(12), ocupation_ne85 => ocupation(47), ocupation_ne100 => ocupation(41), ocupation_ne101 => ocupation(42), ocupation_ne44 => ocupation(15), ocupation_ne110 => ocupation(52), ocupation_ne26 => ocupation(9), ocupation_ne65 => ocupation(20), ocupation_ne48 => ocupation(17), ocupation_ne43 => ocupation(14), ocupation_ne102 => ocupation(43), correspondence_C100 => state_C100, correspondence_S105 => state_S105, correspondence_C138 => state_C138, correspondence_L29 => state_L29, correspondence_S93 => state_S93, Sw04_state => state_Sw04, Sw05_state => state_Sw05, Sw09_state => state_Sw09, Sw41_state => state_Sw41, s71W01_state => state_71W01, s71W02_state => state_71W02, indication.msb => signals_i.msb(27), indication.lsb => signals_i.lsb(27), command.msb => signals_o.msb(27), command.lsb => signals_o.lsb(27), lock_B130 => B130_locking, correspondence_B130 => state_B130);
	railwaySignal_L28 : railwaySignal_28 port map(clock => clock, reset => reset, R12_command => cmd_R12_L28, ocupation_ne44 => ocupation(15), ocupation_ne101 => ocupation(42), ocupation_ne100 => ocupation(41), correspondence_L40 => state_L40, correspondence_S139 => state_S139, indication.msb => signals_i.msb(28), indication.lsb => signals_i.lsb(28), command.msb => signals_o.msb(28), command.lsb => signals_o.lsb(28), lock_L28 => L28_locking, correspondence_L28 => state_L28);
	railwaySignal_S105 : railwaySignal_29 port map(clock => clock, reset => reset, R61_command => cmd_R61_S105, R62_command => cmd_R62_S105, ocupation_ne44 => ocupation(15), ocupation_ne43 => ocupation(14), ocupation_ne48 => ocupation(17), ocupation_ne102 => ocupation(43), ocupation_ne65 => ocupation(20), ocupation_ne26 => ocupation(9), ocupation_ne23 => ocupation(7), ocupation_ne24 => ocupation(8), correspondence_L29 => state_L29, correspondence_S93 => state_S93, correspondence_B89 => state_B89, correspondence_P63 => state_P63, s71W01_state => state_71W01, s71W02_state => state_71W02, s70W02_state => state_70W02, indication.msb => signals_i.msb(29), indication.lsb => signals_i.lsb(29), command.msb => signals_o.msb(29), command.lsb => signals_o.lsb(29), lock_S105 => S105_locking, correspondence_S105 => state_S105);
	railwaySignal_T11 : railwaySignal_30 port map(clock => clock, reset => reset, ocupation_ne47 => ocupation(16), indication.msb => signals_i.msb(30), indication.lsb => signals_i.lsb(30), command.msb => signals_o.msb(30), command.lsb => signals_o.lsb(30), lock_T11 => T11_locking, correspondence_T11 => state_T11);
	railwaySignal_T12 : railwaySignal_31 port map(clock => clock, reset => reset, R4_command => cmd_R4_T12, ocupation_ne47 => ocupation(16), ocupation_ne48 => ocupation(17), correspondence_L29 => state_L29, s71W02_state => state_71W02, indication.msb => signals_i.msb(31), indication.lsb => signals_i.lsb(31), command.msb => signals_o.msb(31), command.lsb => signals_o.lsb(31), lock_T12 => T12_locking, correspondence_T12 => state_T12);
	railwaySignal_L29 : railwaySignal_32 port map(clock => clock, reset => reset, ocupation_ne48 => ocupation(17), indication.msb => signals_i.msb(32), indication.lsb => signals_i.lsb(32), command.msb => signals_o.msb(32), command.lsb => signals_o.lsb(32), lock_L29 => L29_locking, correspondence_L29 => state_L29);
	railwaySignal_S83 : railwaySignal_33 port map(clock => clock, reset => reset, R42_command => cmd_R42_S83, R43_command => cmd_R43_S83, ocupation_ne59 => ocupation(18), ocupation_ne11 => ocupation(4), ocupation_ne52 => ocupation(50), ocupation_ne17 => ocupation(6), ocupation_ne77 => ocupation(48), ocupation_ne78 => ocupation(23), correspondence_S146 => state_S146, correspondence_C109 => state_C109, correspondence_B145 => state_B145, correspondence_L33 => state_L33, s69W03_state => state_69W03, s69W04_state => state_69W04, Sw03_state => state_Sw03, Sw06_state => state_Sw06, indication.msb => signals_i.msb(33), indication.lsb => signals_i.lsb(33), command.msb => signals_o.msb(33), command.lsb => signals_o.lsb(33), lock_S83 => S83_locking, correspondence_S83 => state_S83);
	railwaySignal_S90 : railwaySignal_34 port map(clock => clock, reset => reset, R47_command => cmd_R47_S90, R48_command => cmd_R48_S90, ocupation_ne64 => ocupation(19), ocupation_ne23 => ocupation(7), ocupation_ne24 => ocupation(8), ocupation_ne26 => ocupation(9), correspondence_P60 => state_P60, correspondence_B92 => state_B92, correspondence_L27 => state_L27, s70W01_state => state_70W01, s70W02_state => state_70W02, indication.msb => signals_i.msb(34), indication.lsb => signals_i.lsb(34), command.msb => signals_o.msb(34), command.lsb => signals_o.lsb(34), lock_S90 => S90_locking, correspondence_S90 => state_S90);
	railwaySignal_L30 : railwaySignal_35 port map(clock => clock, reset => reset, R13_command => cmd_R13_L30, ocupation_ne65 => ocupation(20), ocupation_ne102 => ocupation(43), ocupation_ne44 => ocupation(15), correspondence_C104 => state_C104, correspondence_L28 => state_L28, s71W01_state => state_71W01, indication.msb => signals_i.msb(35), indication.lsb => signals_i.lsb(35), command.msb => signals_o.msb(35), command.lsb => signals_o.lsb(35), lock_L30 => L30_locking, correspondence_L30 => state_L30);
	railwaySignal_P64 : railwaySignal_36 port map(clock => clock, reset => reset, R29_command => cmd_R29_P64, ocupation_ne67 => ocupation(21), ocupation_ne70 => ocupation(22), ocupation_ne104 => ocupation(49), ocupation_ne21 => ocupation(51), correspondence_L32 => state_L32, correspondence_P73 => state_P73, Sw03_state => state_Sw03, indication.msb => signals_i.msb(36), indication.lsb => signals_i.lsb(36), command.msb => signals_o.msb(36), command.lsb => signals_o.lsb(36), lock_P64 => P64_locking, correspondence_P64 => state_P64);
	railwaySignal_P65 : railwaySignal_37 port map(clock => clock, reset => reset, R30_command => cmd_R30_P65, ocupation_ne67 => ocupation(21), ocupation_ne103 => ocupation(44), ocupation_ne64 => ocupation(19), correspondence_L41 => state_L41, correspondence_S90 => state_S90, indication.msb => signals_i.msb(37), indication.lsb => signals_i.lsb(37), command.msb => signals_o.msb(37), command.lsb => signals_o.lsb(37), lock_P65 => P65_locking, correspondence_P65 => state_P65);
	railwaySignal_L32 : railwaySignal_38 port map(clock => clock, reset => reset, R14_command => cmd_R14_L32, ocupation_ne70 => ocupation(22), ocupation_ne104 => ocupation(49), ocupation_ne21 => ocupation(51), ocupation_ne94 => ocupation(35), ocupation_ne79 => ocupation(24), ocupation_ne78 => ocupation(23), ocupation_ne99 => ocupation(40), ocupation_ne97 => ocupation(38), correspondence_P73 => state_P73, correspondence_L33 => state_L33, correspondence_P69 => state_P69, Sw03_state => state_Sw03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication.msb => signals_i.msb(38), indication.lsb => signals_i.lsb(38), command.msb => signals_o.msb(38), command.lsb => signals_o.lsb(38), lock_L32 => L32_locking, correspondence_L32 => state_L32);
	railwaySignal_L33 : railwaySignal_39 port map(clock => clock, reset => reset, R15_command => cmd_R15_L33, ocupation_ne78 => ocupation(23), ocupation_ne93 => ocupation(34), ocupation_ne96 => ocupation(37), correspondence_L34 => state_L34, correspondence_P71 => state_P71, indication.msb => signals_i.msb(39), indication.lsb => signals_i.lsb(39), command.msb => signals_o.msb(39), command.lsb => signals_o.lsb(39), lock_L33 => L33_locking, correspondence_L33 => state_L33);
	railwaySignal_S110 : railwaySignal_40 port map(clock => clock, reset => reset, R64_command => cmd_R64_S110, R65_command => cmd_R65_S110, R66_command => cmd_R66_S110, ocupation_ne78 => ocupation(23), ocupation_ne17 => ocupation(6), ocupation_ne79 => ocupation(24), ocupation_ne77 => ocupation(48), ocupation_ne21 => ocupation(51), ocupation_ne95 => ocupation(36), ocupation_ne59 => ocupation(18), ocupation_ne52 => ocupation(50), correspondence_C82 => state_C82, correspondence_B133 => state_B133, correspondence_P72 => state_P72, correspondence_X51 => state_X51, correspondence_S86 => state_S86, correspondence_S144 => state_S144, Sw06_state => state_Sw06, s69W03_state => state_69W03, Sw07_state => state_Sw07, Sw03_state => state_Sw03, indication.msb => signals_i.msb(40), indication.lsb => signals_i.lsb(40), command.msb => signals_o.msb(40), command.lsb => signals_o.lsb(40), lock_S110 => S110_locking, correspondence_S110 => state_S110);
	railwaySignal_C95 : railwaySignal_41 port map(clock => clock, reset => reset, R52_command => cmd_R52_C95, ocupation_ne83 => ocupation(26), ocupation_ne30 => ocupation(11), ocupation_ne90 => ocupation(32), ocupation_ne91 => ocupation(33), ocupation_ne86 => ocupation(28), ocupation_ne87 => ocupation(29), ocupation_ne89 => ocupation(31), correspondence_S122 => state_S122, correspondence_T19 => state_T19, correspondence_T15 => state_T15, correspondence_T21 => state_T21, Sw08_state => state_Sw08, Sw12_state => state_Sw12, Sw11_state => state_Sw11, Sw13_state => state_Sw13, indication.msb => signals_i.msb(41), indication.lsb => signals_i.lsb(41), command.msb => signals_o.msb(41), command.lsb => signals_o.lsb(41), lock_C95 => C95_locking, correspondence_C95 => state_C95);
	railwaySignal_C114 : railwaySignal_42 port map(clock => clock, reset => reset, R67_command => cmd_R67_C114, ocupation_ne83 => ocupation(26), ocupation_ne32 => ocupation(12), ocupation_ne110 => ocupation(52), correspondence_C100 => state_C100, correspondence_C138 => state_C138, Sw04_state => state_Sw04, Sw09_state => state_Sw09, indication.msb => signals_i.msb(42), indication.lsb => signals_i.lsb(42), command.msb => signals_o.msb(42), command.lsb => signals_o.lsb(42), lock_C114 => C114_locking, correspondence_C114 => state_C114);
	railwaySignal_T13 : railwaySignal_43 port map(clock => clock, reset => reset, ocupation_ne84 => ocupation(27), indication.msb => signals_i.msb(43), indication.lsb => signals_i.lsb(43), command.msb => signals_o.msb(43), command.lsb => signals_o.lsb(43), lock_T13 => T13_locking, correspondence_T13 => state_T13);
	railwaySignal_T14 : railwaySignal_44 port map(clock => clock, reset => reset, R5_command => cmd_R5_T14, R6_command => cmd_R6_T14, ocupation_ne84 => ocupation(27), ocupation_ne82 => ocupation(25), ocupation_ne32 => ocupation(12), ocupation_ne85 => ocupation(47), ocupation_ne100 => ocupation(41), ocupation_ne101 => ocupation(42), ocupation_ne44 => ocupation(15), ocupation_ne110 => ocupation(52), ocupation_ne26 => ocupation(9), ocupation_ne65 => ocupation(20), ocupation_ne48 => ocupation(17), ocupation_ne43 => ocupation(14), ocupation_ne102 => ocupation(43), correspondence_C100 => state_C100, correspondence_S105 => state_S105, correspondence_C138 => state_C138, correspondence_L29 => state_L29, correspondence_S93 => state_S93, Sw04_state => state_Sw04, Sw05_state => state_Sw05, Sw09_state => state_Sw09, Sw41_state => state_Sw41, s71W01_state => state_71W01, s71W02_state => state_71W02, indication.msb => signals_i.msb(44), indication.lsb => signals_i.lsb(44), command.msb => signals_o.msb(44), command.lsb => signals_o.lsb(44), lock_T14 => T14_locking, correspondence_T14 => state_T14);
	railwaySignal_T15 : railwaySignal_45 port map(clock => clock, reset => reset, ocupation_ne86 => ocupation(28), indication.msb => signals_i.msb(45), indication.lsb => signals_i.lsb(45), command.msb => signals_o.msb(45), command.lsb => signals_o.lsb(45), lock_T15 => T15_locking, correspondence_T15 => state_T15);
	railwaySignal_S119 : railwaySignal_46 port map(clock => clock, reset => reset, R72_command => cmd_R72_S119, R73_command => cmd_R73_S119, ocupation_ne86 => ocupation(28), ocupation_ne88 => ocupation(30), ocupation_ne87 => ocupation(29), ocupation_ne91 => ocupation(33), ocupation_ne30 => ocupation(11), ocupation_ne29 => ocupation(10), ocupation_ne110 => ocupation(52), ocupation_ne83 => ocupation(26), correspondence_T17 => state_T17, correspondence_S97 => state_S97, correspondence_C138 => state_C138, correspondence_C114 => state_C114, Sw11_state => state_Sw11, Sw12_state => state_Sw12, Sw13_state => state_Sw13, Sw08_state => state_Sw08, Sw09_state => state_Sw09, indication.msb => signals_i.msb(46), indication.lsb => signals_i.lsb(46), command.msb => signals_o.msb(46), command.lsb => signals_o.lsb(46), lock_S119 => S119_locking, correspondence_S119 => state_S119);
	railwaySignal_T17 : railwaySignal_47 port map(clock => clock, reset => reset, ocupation_ne88 => ocupation(30), indication.msb => signals_i.msb(47), indication.lsb => signals_i.lsb(47), command.msb => signals_o.msb(47), command.lsb => signals_o.lsb(47), lock_T17 => T17_locking, correspondence_T17 => state_T17);
	railwaySignal_C118 : railwaySignal_48 port map(clock => clock, reset => reset, R71_command => cmd_R71_C118, ocupation_ne88 => ocupation(30), ocupation_ne86 => ocupation(28), correspondence_T15 => state_T15, Sw11_state => state_Sw11, indication.msb => signals_i.msb(48), indication.lsb => signals_i.lsb(48), command.msb => signals_o.msb(48), command.lsb => signals_o.lsb(48), lock_C118 => C118_locking, correspondence_C118 => state_C118);
	railwaySignal_T19 : railwaySignal_49 port map(clock => clock, reset => reset, ocupation_ne89 => ocupation(31), indication.msb => signals_i.msb(49), indication.lsb => signals_i.lsb(49), command.msb => signals_o.msb(49), command.lsb => signals_o.lsb(49), lock_T19 => T19_locking, correspondence_T19 => state_T19);
	railwaySignal_T20 : railwaySignal_50 port map(clock => clock, reset => reset, R7_command => cmd_R7_T20, ocupation_ne89 => ocupation(31), ocupation_ne30 => ocupation(11), ocupation_ne29 => ocupation(10), ocupation_ne110 => ocupation(52), ocupation_ne83 => ocupation(26), correspondence_S97 => state_S97, correspondence_C138 => state_C138, correspondence_C114 => state_C114, Sw12_state => state_Sw12, Sw08_state => state_Sw08, Sw09_state => state_Sw09, indication.msb => signals_i.msb(50), indication.lsb => signals_i.lsb(50), command.msb => signals_o.msb(50), command.lsb => signals_o.lsb(50), lock_T20 => T20_locking, correspondence_T20 => state_T20);
	railwaySignal_T21 : railwaySignal_51 port map(clock => clock, reset => reset, ocupation_ne90 => ocupation(32), indication.msb => signals_i.msb(51), indication.lsb => signals_i.lsb(51), command.msb => signals_o.msb(51), command.lsb => signals_o.lsb(51), lock_T21 => T21_locking, correspondence_T21 => state_T21);
	railwaySignal_T22 : railwaySignal_52 port map(clock => clock, reset => reset, R8_command => cmd_R8_T22, ocupation_ne90 => ocupation(32), ocupation_ne91 => ocupation(33), ocupation_ne30 => ocupation(11), ocupation_ne29 => ocupation(10), ocupation_ne110 => ocupation(52), ocupation_ne83 => ocupation(26), correspondence_S97 => state_S97, correspondence_C138 => state_C138, correspondence_C114 => state_C114, Sw12_state => state_Sw12, Sw13_state => state_Sw13, Sw08_state => state_Sw08, Sw09_state => state_Sw09, indication.msb => signals_i.msb(52), indication.lsb => signals_i.lsb(52), command.msb => signals_o.msb(52), command.lsb => signals_o.lsb(52), lock_T22 => T22_locking, correspondence_T22 => state_T22);
	railwaySignal_L34 : railwaySignal_53 port map(clock => clock, reset => reset, R16_command => cmd_R16_L34, ocupation_ne93 => ocupation(34), ocupation_ne96 => ocupation(37), ocupation_ne98 => ocupation(39), correspondence_P71 => state_P71, correspondence_L38 => state_L38, indication.msb => signals_i.msb(53), indication.lsb => signals_i.lsb(53), command.msb => signals_o.msb(53), command.lsb => signals_o.lsb(53), lock_L34 => L34_locking, correspondence_L34 => state_L34);
	railwaySignal_S135 : railwaySignal_54 port map(clock => clock, reset => reset, R82_command => cmd_R82_S135, R83_command => cmd_R83_S135, ocupation_ne94 => ocupation(35), ocupation_ne77 => ocupation(48), ocupation_ne21 => ocupation(51), ocupation_ne52 => ocupation(50), correspondence_B133 => state_B133, correspondence_P72 => state_P72, correspondence_S86 => state_S86, correspondence_S144 => state_S144, Sw07_state => state_Sw07, Sw03_state => state_Sw03, indication.msb => signals_i.msb(54), indication.lsb => signals_i.lsb(54), command.msb => signals_o.msb(54), command.lsb => signals_o.lsb(54), lock_S135 => S135_locking, correspondence_S135 => state_S135);
	railwaySignal_L35 : railwaySignal_55 port map(clock => clock, reset => reset, R17_command => cmd_R17_L35, ocupation_ne95 => ocupation(36), ocupation_ne59 => ocupation(18), correspondence_X50 => state_X50, correspondence_S83 => state_S83, indication.msb => signals_i.msb(55), indication.lsb => signals_i.lsb(55), command.msb => signals_o.msb(55), command.lsb => signals_o.lsb(55), lock_L35 => L35_locking, correspondence_L35 => state_L35);
	railwaySignal_X50 : railwaySignal_56 port map(clock => clock, reset => reset, R25_command => cmd_R25_X50, ocupation_ne95 => ocupation(36), ocupation_ne59 => ocupation(18), ocupation_ne11 => ocupation(4), ocupation_ne17 => ocupation(6), ocupation_ne52 => ocupation(50), correspondence_S83 => state_S83, correspondence_S146 => state_S146, correspondence_C109 => state_C109, s69W03_state => state_69W03, s69W04_state => state_69W04, Lc01_state => state_Lc01, indication.msb => signals_i.msb(56), indication.lsb => signals_i.lsb(56), command.msb => signals_o.msb(56), command.lsb => signals_o.lsb(56), lock_X50 => X50_locking, correspondence_X50 => state_X50);
	railwaySignal_X51 : railwaySignal_57 port map(clock => clock, reset => reset, R26_command => cmd_R26_X51, ocupation_ne95 => ocupation(36), ocupation_ne9 => ocupation(3), ocupation_ne1 => ocupation(0), ocupation_ne7 => ocupation(2), correspondence_S80 => state_S80, correspondence_T01 => state_T01, correspondence_T05 => state_T05, s68W02_state => state_68W02, Lc01_state => state_Lc01, indication.msb => signals_i.msb(57), indication.lsb => signals_i.lsb(57), command.msb => signals_o.msb(57), command.lsb => signals_o.lsb(57), lock_X51 => X51_locking, correspondence_X51 => state_X51);
	railwaySignal_P70 : railwaySignal_58 port map(clock => clock, reset => reset, R33_command => cmd_R33_P70, ocupation_ne96 => ocupation(37), ocupation_ne93 => ocupation(34), ocupation_ne78 => ocupation(23), ocupation_ne79 => ocupation(24), ocupation_ne21 => ocupation(51), ocupation_ne17 => ocupation(6), ocupation_ne77 => ocupation(48), correspondence_S110 => state_S110, correspondence_C82 => state_C82, correspondence_B133 => state_B133, correspondence_P72 => state_P72, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication.msb => signals_i.msb(58), indication.lsb => signals_i.lsb(58), command.msb => signals_o.msb(58), command.lsb => signals_o.lsb(58), lock_P70 => P70_locking, correspondence_P70 => state_P70);
	railwaySignal_P71 : railwaySignal_59 port map(clock => clock, reset => reset, R34_command => cmd_R34_P71, ocupation_ne96 => ocupation(37), ocupation_ne98 => ocupation(39), ocupation_ne105 => ocupation(45), correspondence_L38 => state_L38, correspondence_T23 => state_T23, indication.msb => signals_i.msb(59), indication.lsb => signals_i.lsb(59), command.msb => signals_o.msb(59), command.lsb => signals_o.lsb(59), lock_P71 => P71_locking, correspondence_P71 => state_P71);
	railwaySignal_L37 : railwaySignal_60 port map(clock => clock, reset => reset, R18_command => cmd_R18_L37, ocupation_ne97 => ocupation(38), ocupation_ne94 => ocupation(35), ocupation_ne21 => ocupation(51), ocupation_ne77 => ocupation(48), correspondence_S135 => state_S135, correspondence_B133 => state_B133, correspondence_P72 => state_P72, Sw07_state => state_Sw07, indication.msb => signals_i.msb(60), indication.lsb => signals_i.lsb(60), command.msb => signals_o.msb(60), command.lsb => signals_o.lsb(60), lock_L37 => L37_locking, correspondence_L37 => state_L37);
	railwaySignal_L38 : railwaySignal_61 port map(clock => clock, reset => reset, R19_command => cmd_R19_L38, ocupation_ne98 => ocupation(39), ocupation_ne105 => ocupation(45), correspondence_T23 => state_T23, indication.msb => signals_i.msb(61), indication.lsb => signals_i.lsb(61), command.msb => signals_o.msb(61), command.lsb => signals_o.lsb(61), lock_L38 => L38_locking, correspondence_L38 => state_L38);
	railwaySignal_P68 : railwaySignal_62 port map(clock => clock, reset => reset, R31_command => cmd_R31_P68, ocupation_ne99 => ocupation(40), ocupation_ne97 => ocupation(38), ocupation_ne94 => ocupation(35), correspondence_L37 => state_L37, correspondence_S135 => state_S135, indication.msb => signals_i.msb(62), indication.lsb => signals_i.lsb(62), command.msb => signals_o.msb(62), command.lsb => signals_o.lsb(62), lock_P68 => P68_locking, correspondence_P68 => state_P68);
	railwaySignal_P69 : railwaySignal_63 port map(clock => clock, reset => reset, R32_command => cmd_R32_P69, ocupation_ne99 => ocupation(40), ocupation_ne106 => ocupation(46), ocupation_ne4 => ocupation(1), correspondence_T03 => state_T03, indication.msb => signals_i.msb(63), indication.lsb => signals_i.lsb(63), command.msb => signals_o.msb(63), command.lsb => signals_o.lsb(63), lock_P69 => P69_locking, correspondence_P69 => state_P69);
	railwaySignal_S139 : railwaySignal_64 port map(clock => clock, reset => reset, R85_command => cmd_R85_S139, R86_command => cmd_R86_S139, ocupation_ne100 => ocupation(41), ocupation_ne110 => ocupation(52), ocupation_ne85 => ocupation(47), ocupation_ne29 => ocupation(10), ocupation_ne32 => ocupation(12), ocupation_ne41 => ocupation(13), ocupation_ne84 => ocupation(27), correspondence_S102 => state_S102, correspondence_S131 => state_S131, correspondence_S115 => state_S115, correspondence_B101 => state_B101, correspondence_P58 => state_P58, correspondence_T13 => state_T13, Sw41_state => state_Sw41, Sw09_state => state_Sw09, Sw05_state => state_Sw05, indication.msb => signals_i.msb(64), indication.lsb => signals_i.lsb(64), command.msb => signals_o.msb(64), command.lsb => signals_o.lsb(64), lock_S139 => S139_locking, correspondence_S139 => state_S139);
	railwaySignal_L40 : railwaySignal_65 port map(clock => clock, reset => reset, R20_command => cmd_R20_L40, ocupation_ne101 => ocupation(42), ocupation_ne100 => ocupation(41), ocupation_ne110 => ocupation(52), ocupation_ne85 => ocupation(47), correspondence_S139 => state_S139, correspondence_S102 => state_S102, correspondence_S131 => state_S131, Sw41_state => state_Sw41, indication.msb => signals_i.msb(65), indication.lsb => signals_i.lsb(65), command.msb => signals_o.msb(65), command.lsb => signals_o.lsb(65), lock_L40 => L40_locking, correspondence_L40 => state_L40);
	railwaySignal_C104 : railwaySignal_66 port map(clock => clock, reset => reset, R60_command => cmd_R60_C104, ocupation_ne102 => ocupation(43), ocupation_ne44 => ocupation(15), ocupation_ne101 => ocupation(42), correspondence_L28 => state_L28, correspondence_L40 => state_L40, s71W01_state => state_71W01, indication.msb => signals_i.msb(66), indication.lsb => signals_i.lsb(66), command.msb => signals_o.msb(66), command.lsb => signals_o.lsb(66), lock_C104 => C104_locking, correspondence_C104 => state_C104);
	railwaySignal_L41 : railwaySignal_67 port map(clock => clock, reset => reset, R21_command => cmd_R21_L41, ocupation_ne103 => ocupation(44), ocupation_ne64 => ocupation(19), ocupation_ne23 => ocupation(7), ocupation_ne24 => ocupation(8), correspondence_S90 => state_S90, correspondence_P60 => state_P60, correspondence_B92 => state_B92, s70W01_state => state_70W01, indication.msb => signals_i.msb(67), indication.lsb => signals_i.lsb(67), command.msb => signals_o.msb(67), command.lsb => signals_o.lsb(67), lock_L41 => L41_locking, correspondence_L41 => state_L41);
	railwaySignal_T23 : railwaySignal_68 port map(clock => clock, reset => reset, ocupation_ne105 => ocupation(45), indication.msb => signals_i.msb(68), indication.lsb => signals_i.lsb(68), command.msb => signals_o.msb(68), command.lsb => signals_o.lsb(68), lock_T23 => T23_locking, correspondence_T23 => state_T23);
	railwaySignal_T24 : railwaySignal_69 port map(clock => clock, reset => reset, R9_command => cmd_R9_T24, ocupation_ne105 => ocupation(45), ocupation_ne98 => ocupation(39), ocupation_ne96 => ocupation(37), ocupation_ne78 => ocupation(23), ocupation_ne93 => ocupation(34), correspondence_P70 => state_P70, correspondence_S110 => state_S110, indication.msb => signals_i.msb(69), indication.lsb => signals_i.lsb(69), command.msb => signals_o.msb(69), command.lsb => signals_o.lsb(69), lock_T24 => T24_locking, correspondence_T24 => state_T24);
	railwaySignal_L42 : railwaySignal_70 port map(clock => clock, reset => reset, R22_command => cmd_R22_L42, ocupation_ne106 => ocupation(46), ocupation_ne99 => ocupation(40), ocupation_ne97 => ocupation(38), correspondence_P68 => state_P68, correspondence_L37 => state_L37, indication.msb => signals_i.msb(70), indication.lsb => signals_i.lsb(70), command.msb => signals_o.msb(70), command.lsb => signals_o.lsb(70), lock_L42 => L42_locking, correspondence_L42 => state_L42);
	railwaySignal_S131 : railwaySignal_71 port map(clock => clock, reset => reset, R79_command => cmd_R79_S131, R80_command => cmd_R80_S131, ocupation_ne85 => ocupation(47), ocupation_ne41 => ocupation(13), ocupation_ne84 => ocupation(27), correspondence_P58 => state_P58, correspondence_T13 => state_T13, Sw05_state => state_Sw05, indication.msb => signals_i.msb(71), indication.lsb => signals_i.lsb(71), command.msb => signals_o.msb(71), command.lsb => signals_o.lsb(71), lock_S131 => S131_locking, correspondence_S131 => state_S131);
	railwaySignal_B133 : railwaySignal_72 port map(clock => clock, reset => reset, R81_command => cmd_R81_B133, ocupation_ne77 => ocupation(48), ocupation_ne52 => ocupation(50), ocupation_ne95 => ocupation(36), ocupation_ne11 => ocupation(4), ocupation_ne14 => ocupation(5), ocupation_ne59 => ocupation(18), correspondence_S86 => state_S86, correspondence_X51 => state_X51, correspondence_T07 => state_T07, Sw03_state => state_Sw03, s69W03_state => state_69W03, s69W04_state => state_69W04, indication.msb => signals_i.msb(72), indication.lsb => signals_i.lsb(72), command.msb => signals_o.msb(72), command.lsb => signals_o.lsb(72), lock_B133 => B133_locking, correspondence_B133 => state_B133);
	railwaySignal_B145 : railwaySignal_73 port map(clock => clock, reset => reset, R89_command => cmd_R89_B145, R90_command => cmd_R90_B145, ocupation_ne77 => ocupation(48), ocupation_ne79 => ocupation(24), ocupation_ne78 => ocupation(23), ocupation_ne94 => ocupation(35), ocupation_ne97 => ocupation(38), ocupation_ne99 => ocupation(40), ocupation_ne93 => ocupation(34), ocupation_ne4 => ocupation(1), ocupation_ne106 => ocupation(46), correspondence_L33 => state_L33, correspondence_P69 => state_P69, correspondence_L34 => state_L34, correspondence_T03 => state_T03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication.msb => signals_i.msb(73), indication.lsb => signals_i.lsb(73), command.msb => signals_o.msb(73), command.lsb => signals_o.lsb(73), lock_B145 => B145_locking, correspondence_B145 => state_B145);
	railwaySignal_B143 : railwaySignal_74 port map(clock => clock, reset => reset, R87_command => cmd_R87_B143, ocupation_ne104 => ocupation(49), ocupation_ne70 => ocupation(22), ocupation_ne21 => ocupation(51), correspondence_L32 => state_L32, correspondence_P73 => state_P73, Sw03_state => state_Sw03, indication.msb => signals_i.msb(74), indication.lsb => signals_i.lsb(74), command.msb => signals_o.msb(74), command.lsb => signals_o.lsb(74), lock_B143 => B143_locking, correspondence_B143 => state_B143);
	railwaySignal_S86 : railwaySignal_75 port map(clock => clock, reset => reset, R44_command => cmd_R44_S86, R45_command => cmd_R45_S86, ocupation_ne52 => ocupation(50), ocupation_ne11 => ocupation(4), ocupation_ne59 => ocupation(18), ocupation_ne95 => ocupation(36), ocupation_ne14 => ocupation(5), ocupation_ne9 => ocupation(3), correspondence_X51 => state_X51, correspondence_T07 => state_T07, correspondence_S80 => state_S80, s69W03_state => state_69W03, s69W04_state => state_69W04, Lc01_state => state_Lc01, indication.msb => signals_i.msb(75), indication.lsb => signals_i.lsb(75), command.msb => signals_o.msb(75), command.lsb => signals_o.lsb(75), lock_S86 => S86_locking, correspondence_S86 => state_S86);
	railwaySignal_S146 : railwaySignal_76 port map(clock => clock, reset => reset, R91_command => cmd_R91_S146, ocupation_ne52 => ocupation(50), ocupation_ne77 => ocupation(48), ocupation_ne94 => ocupation(35), ocupation_ne79 => ocupation(24), ocupation_ne78 => ocupation(23), ocupation_ne99 => ocupation(40), ocupation_ne97 => ocupation(38), correspondence_B145 => state_B145, correspondence_L33 => state_L33, correspondence_P69 => state_P69, Sw03_state => state_Sw03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication.msb => signals_i.msb(76), indication.lsb => signals_i.lsb(76), command.msb => signals_o.msb(76), command.lsb => signals_o.lsb(76), lock_S146 => S146_locking, correspondence_S146 => state_S146);
	railwaySignal_P72 : railwaySignal_77 port map(clock => clock, reset => reset, R35_command => cmd_R35_P72, ocupation_ne21 => ocupation(51), ocupation_ne104 => ocupation(49), correspondence_S144 => state_S144, correspondence_B143 => state_B143, Sw03_state => state_Sw03, indication.msb => signals_i.msb(77), indication.lsb => signals_i.lsb(77), command.msb => signals_o.msb(77), command.lsb => signals_o.lsb(77), lock_P72 => P72_locking, correspondence_P72 => state_P72);
	railwaySignal_P73 : railwaySignal_78 port map(clock => clock, reset => reset, R36_command => cmd_R36_P73, R37_command => cmd_R37_P73, ocupation_ne21 => ocupation(51), ocupation_ne79 => ocupation(24), ocupation_ne78 => ocupation(23), ocupation_ne94 => ocupation(35), ocupation_ne97 => ocupation(38), ocupation_ne99 => ocupation(40), ocupation_ne93 => ocupation(34), ocupation_ne4 => ocupation(1), ocupation_ne106 => ocupation(46), correspondence_L33 => state_L33, correspondence_P69 => state_P69, correspondence_L34 => state_L34, correspondence_T03 => state_T03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication.msb => signals_i.msb(78), indication.lsb => signals_i.lsb(78), command.msb => signals_o.msb(78), command.lsb => signals_o.lsb(78), lock_P73 => P73_locking, correspondence_P73 => state_P73);
	railwaySignal_S144 : railwaySignal_79 port map(clock => clock, reset => reset, R88_command => cmd_R88_S144, ocupation_ne21 => ocupation(51), ocupation_ne104 => ocupation(49), ocupation_ne70 => ocupation(22), correspondence_B143 => state_B143, correspondence_L32 => state_L32, Sw03_state => state_Sw03, indication.msb => signals_i.msb(79), indication.lsb => signals_i.lsb(79), command.msb => signals_o.msb(79), command.lsb => signals_o.lsb(79), lock_S144 => S144_locking, correspondence_S144 => state_S144);
	railwaySignal_S102 : railwaySignal_80 port map(clock => clock, reset => reset, R58_command => cmd_R58_S102, R59_command => cmd_R59_S102, ocupation_ne110 => ocupation(52), ocupation_ne32 => ocupation(12), ocupation_ne29 => ocupation(10), ocupation_ne82 => ocupation(25), ocupation_ne41 => ocupation(13), ocupation_ne83 => ocupation(26), ocupation_ne84 => ocupation(27), correspondence_S115 => state_S115, correspondence_B101 => state_B101, correspondence_C95 => state_C95, correspondence_P58 => state_P58, correspondence_T13 => state_T13, correspondence_B96 => state_B96, Sw09_state => state_Sw09, Sw04_state => state_Sw04, Sw05_state => state_Sw05, indication.msb => signals_i.msb(80), indication.lsb => signals_i.lsb(80), command.msb => signals_o.msb(80), command.lsb => signals_o.lsb(80), lock_S102 => S102_locking, correspondence_S102 => state_S102);
	railwaySignal_C138 : railwaySignal_81 port map(clock => clock, reset => reset, R84_command => cmd_R84_C138, ocupation_ne110 => ocupation(52), ocupation_ne100 => ocupation(41), ocupation_ne101 => ocupation(42), ocupation_ne44 => ocupation(15), ocupation_ne26 => ocupation(9), ocupation_ne65 => ocupation(20), ocupation_ne48 => ocupation(17), ocupation_ne43 => ocupation(14), ocupation_ne102 => ocupation(43), correspondence_S105 => state_S105, correspondence_L29 => state_L29, correspondence_S93 => state_S93, Sw41_state => state_Sw41, s71W01_state => state_71W01, s71W02_state => state_71W02, indication.msb => signals_i.msb(81), indication.lsb => signals_i.lsb(81), command.msb => signals_o.msb(81), command.lsb => signals_o.lsb(81), lock_C138 => C138_locking, correspondence_C138 => state_C138);
	node_ne1 : node_0 port map(clock => clock, ocupation => ocupation(0), reset => reset, R1_command => cmd_R1_ne1, R38_command => cmd_R38_ne1, R39_command => cmd_R39_ne1, state => state_ne1, locking => ne1_locking);
	node_ne4 : node_1 port map(clock => clock, ocupation => ocupation(1), reset => reset, R10_command => cmd_R10_ne4, R32_command => cmd_R32_ne4, state => state_ne4, locking => ne4_locking);
	node_ne7 : node_2 port map(clock => clock, ocupation => ocupation(2), reset => reset, R2_command => cmd_R2_ne7, R23_command => cmd_R23_ne7, R40_command => cmd_R40_ne7, state => state_ne7, locking => ne7_locking);
	node_ne9 : node_3 port map(clock => clock, ocupation => ocupation(3), reset => reset, R23_command => cmd_R23_ne9, R24_command => cmd_R24_ne9, R26_command => cmd_R26_ne9, R38_command => cmd_R38_ne9, R39_command => cmd_R39_ne9, R40_command => cmd_R40_ne9, state => state_ne9, locking => ne9_locking);
	node_ne11 : node_4 port map(clock => clock, ocupation => ocupation(4), reset => reset, R42_command => cmd_R42_ne11, R44_command => cmd_R44_ne11, state => state_ne11, locking => ne11_locking);
	node_ne14 : node_5 port map(clock => clock, ocupation => ocupation(5), reset => reset, R3_command => cmd_R3_ne14, R45_command => cmd_R45_ne14, state => state_ne14, locking => ne14_locking);
	node_ne17 : node_6 port map(clock => clock, ocupation => ocupation(6), reset => reset, R41_command => cmd_R41_ne17, R43_command => cmd_R43_ne17, R63_command => cmd_R63_ne17, R64_command => cmd_R64_ne17, state => state_ne17, locking => ne17_locking);
	node_ne23 : node_7 port map(clock => clock, ocupation => ocupation(7), reset => reset, R27_command => cmd_R27_ne23, R46_command => cmd_R46_ne23, R47_command => cmd_R47_ne23, R50_command => cmd_R50_ne23, state => state_ne23, locking => ne23_locking);
	node_ne24 : node_8 port map(clock => clock, ocupation => ocupation(8), reset => reset, R28_command => cmd_R28_ne24, R48_command => cmd_R48_ne24, R49_command => cmd_R49_ne24, R51_command => cmd_R51_ne24, state => state_ne24, locking => ne24_locking);
	node_ne26 : node_9 port map(clock => clock, ocupation => ocupation(9), reset => reset, R11_command => cmd_R11_ne26, R27_command => cmd_R27_ne26, R49_command => cmd_R49_ne26, R50_command => cmd_R50_ne26, R51_command => cmd_R51_ne26, R62_command => cmd_R62_ne26, state => state_ne26, locking => ne26_locking);
	node_ne29 : node_10 port map(clock => clock, ocupation => ocupation(10), reset => reset, R53_command => cmd_R53_ne29, R54_command => cmd_R54_ne29, R57_command => cmd_R57_ne29, R59_command => cmd_R59_ne29, state => state_ne29, locking => ne29_locking);
	node_ne30 : node_11 port map(clock => clock, ocupation => ocupation(11), reset => reset, R7_command => cmd_R7_ne30, R8_command => cmd_R8_ne30, R52_command => cmd_R52_ne30, R53_command => cmd_R53_ne30, R54_command => cmd_R54_ne30, R55_command => cmd_R55_ne30, R73_command => cmd_R73_ne30, R74_command => cmd_R74_ne30, R75_command => cmd_R75_ne30, R76_command => cmd_R76_ne30, state => state_ne30, locking => ne30_locking);
	node_ne32 : node_12 port map(clock => clock, ocupation => ocupation(12), reset => reset, R5_command => cmd_R5_ne32, R56_command => cmd_R56_ne32, R58_command => cmd_R58_ne32, R67_command => cmd_R67_ne32, R68_command => cmd_R68_ne32, R69_command => cmd_R69_ne32, R70_command => cmd_R70_ne32, R77_command => cmd_R77_ne32, state => state_ne32, locking => ne32_locking);
	node_ne41 : node_13 port map(clock => clock, ocupation => ocupation(13), reset => reset, R69_command => cmd_R69_ne41, R77_command => cmd_R77_ne41, R78_command => cmd_R78_ne41, R79_command => cmd_R79_ne41, state => state_ne41, locking => ne41_locking);
	node_ne43 : node_14 port map(clock => clock, ocupation => ocupation(14), reset => reset, R61_command => cmd_R61_ne43, state => state_ne43, locking => ne43_locking);
	node_ne44 : node_15 port map(clock => clock, ocupation => ocupation(15), reset => reset, R6_command => cmd_R6_ne44, R12_command => cmd_R12_ne44, R60_command => cmd_R60_ne44, R61_command => cmd_R61_ne44, R62_command => cmd_R62_ne44, R78_command => cmd_R78_ne44, R84_command => cmd_R84_ne44, state => state_ne44, locking => ne44_locking);
	node_ne47 : node_16 port map(clock => clock, ocupation => ocupation(16), reset => reset, R4_command => cmd_R4_ne47, state => state_ne47, locking => ne47_locking);
	node_ne48 : node_17 port map(clock => clock, ocupation => ocupation(17), reset => reset, R4_command => cmd_R4_ne48, R61_command => cmd_R61_ne48, state => state_ne48, locking => ne48_locking);
	node_ne59 : node_18 port map(clock => clock, ocupation => ocupation(18), reset => reset, R25_command => cmd_R25_ne59, R41_command => cmd_R41_ne59, R42_command => cmd_R42_ne59, R43_command => cmd_R43_ne59, R44_command => cmd_R44_ne59, state => state_ne59, locking => ne59_locking);
	node_ne64 : node_19 port map(clock => clock, ocupation => ocupation(19), reset => reset, R21_command => cmd_R21_ne64, R28_command => cmd_R28_ne64, R46_command => cmd_R46_ne64, R47_command => cmd_R47_ne64, R48_command => cmd_R48_ne64, state => state_ne64, locking => ne64_locking);
	node_ne65 : node_20 port map(clock => clock, ocupation => ocupation(20), reset => reset, R11_command => cmd_R11_ne65, R13_command => cmd_R13_ne65, R62_command => cmd_R62_ne65, state => state_ne65, locking => ne65_locking);
	node_ne67 : node_21 port map(clock => clock, ocupation => ocupation(21), reset => reset, R28_command => cmd_R28_ne67, R29_command => cmd_R29_ne67, R30_command => cmd_R30_ne67, R46_command => cmd_R46_ne67, state => state_ne67, locking => ne67_locking);
	node_ne70 : node_22 port map(clock => clock, ocupation => ocupation(22), reset => reset, R14_command => cmd_R14_ne70, R29_command => cmd_R29_ne70, R87_command => cmd_R87_ne70, state => state_ne70, locking => ne70_locking);
	node_ne78 : node_23 port map(clock => clock, ocupation => ocupation(23), reset => reset, R15_command => cmd_R15_ne78, R33_command => cmd_R33_ne78, R36_command => cmd_R36_ne78, R63_command => cmd_R63_ne78, R64_command => cmd_R64_ne78, R65_command => cmd_R65_ne78, R66_command => cmd_R66_ne78, R89_command => cmd_R89_ne78, state => state_ne78, locking => ne78_locking);
	node_ne79 : node_24 port map(clock => clock, ocupation => ocupation(24), reset => reset, R36_command => cmd_R36_ne79, R65_command => cmd_R65_ne79, R66_command => cmd_R66_ne79, R89_command => cmd_R89_ne79, state => state_ne79, locking => ne79_locking);
	node_ne82 : node_25 port map(clock => clock, ocupation => ocupation(25), reset => reset, R5_command => cmd_R5_ne82, R69_command => cmd_R69_ne82, R70_command => cmd_R70_ne82, R77_command => cmd_R77_ne82, state => state_ne82, locking => ne82_locking);
	node_ne83 : node_26 port map(clock => clock, ocupation => ocupation(26), reset => reset, R52_command => cmd_R52_ne83, R55_command => cmd_R55_ne83, R67_command => cmd_R67_ne83, R68_command => cmd_R68_ne83, state => state_ne83, locking => ne83_locking);
	node_ne84 : node_27 port map(clock => clock, ocupation => ocupation(27), reset => reset, R5_command => cmd_R5_ne84, R6_command => cmd_R6_ne84, R70_command => cmd_R70_ne84, R80_command => cmd_R80_ne84, state => state_ne84, locking => ne84_locking);
	node_ne86 : node_28 port map(clock => clock, ocupation => ocupation(28), reset => reset, R71_command => cmd_R71_ne86, R72_command => cmd_R72_ne86, R73_command => cmd_R73_ne86, R75_command => cmd_R75_ne86, state => state_ne86, locking => ne86_locking);
	node_ne87 : node_29 port map(clock => clock, ocupation => ocupation(29), reset => reset, R73_command => cmd_R73_ne87, R75_command => cmd_R75_ne87, state => state_ne87, locking => ne87_locking);
	node_ne88 : node_30 port map(clock => clock, ocupation => ocupation(30), reset => reset, R71_command => cmd_R71_ne88, R72_command => cmd_R72_ne88, state => state_ne88, locking => ne88_locking);
	node_ne89 : node_31 port map(clock => clock, ocupation => ocupation(31), reset => reset, R7_command => cmd_R7_ne89, R74_command => cmd_R74_ne89, state => state_ne89, locking => ne89_locking);
	node_ne90 : node_32 port map(clock => clock, ocupation => ocupation(32), reset => reset, R8_command => cmd_R8_ne90, R76_command => cmd_R76_ne90, state => state_ne90, locking => ne90_locking);
	node_ne91 : node_33 port map(clock => clock, ocupation => ocupation(33), reset => reset, R8_command => cmd_R8_ne91, R73_command => cmd_R73_ne91, R75_command => cmd_R75_ne91, R76_command => cmd_R76_ne91, state => state_ne91, locking => ne91_locking);
	node_ne93 : node_34 port map(clock => clock, ocupation => ocupation(34), reset => reset, R15_command => cmd_R15_ne93, R16_command => cmd_R16_ne93, R33_command => cmd_R33_ne93, state => state_ne93, locking => ne93_locking);
	node_ne94 : node_35 port map(clock => clock, ocupation => ocupation(35), reset => reset, R18_command => cmd_R18_ne94, R37_command => cmd_R37_ne94, R82_command => cmd_R82_ne94, R83_command => cmd_R83_ne94, R90_command => cmd_R90_ne94, state => state_ne94, locking => ne94_locking);
	node_ne95 : node_36 port map(clock => clock, ocupation => ocupation(36), reset => reset, R17_command => cmd_R17_ne95, R24_command => cmd_R24_ne95, R25_command => cmd_R25_ne95, R26_command => cmd_R26_ne95, R41_command => cmd_R41_ne95, R44_command => cmd_R44_ne95, state => state_ne95, locking => ne95_locking);
	node_ne96 : node_37 port map(clock => clock, ocupation => ocupation(37), reset => reset, R9_command => cmd_R9_ne96, R16_command => cmd_R16_ne96, R33_command => cmd_R33_ne96, R34_command => cmd_R34_ne96, state => state_ne96, locking => ne96_locking);
	node_ne97 : node_38 port map(clock => clock, ocupation => ocupation(38), reset => reset, R18_command => cmd_R18_ne97, R31_command => cmd_R31_ne97, R37_command => cmd_R37_ne97, R90_command => cmd_R90_ne97, state => state_ne97, locking => ne97_locking);
	node_ne98 : node_39 port map(clock => clock, ocupation => ocupation(39), reset => reset, R9_command => cmd_R9_ne98, R19_command => cmd_R19_ne98, R34_command => cmd_R34_ne98, state => state_ne98, locking => ne98_locking);
	node_ne99 : node_40 port map(clock => clock, ocupation => ocupation(40), reset => reset, R22_command => cmd_R22_ne99, R31_command => cmd_R31_ne99, R32_command => cmd_R32_ne99, R37_command => cmd_R37_ne99, R90_command => cmd_R90_ne99, state => state_ne99, locking => ne99_locking);
	node_ne100 : node_41 port map(clock => clock, ocupation => ocupation(41), reset => reset, R6_command => cmd_R6_ne100, R20_command => cmd_R20_ne100, R78_command => cmd_R78_ne100, R84_command => cmd_R84_ne100, R85_command => cmd_R85_ne100, R86_command => cmd_R86_ne100, state => state_ne100, locking => ne100_locking);
	node_ne101 : node_42 port map(clock => clock, ocupation => ocupation(42), reset => reset, R6_command => cmd_R6_ne101, R12_command => cmd_R12_ne101, R20_command => cmd_R20_ne101, R78_command => cmd_R78_ne101, R84_command => cmd_R84_ne101, state => state_ne101, locking => ne101_locking);
	node_ne102 : node_43 port map(clock => clock, ocupation => ocupation(43), reset => reset, R13_command => cmd_R13_ne102, R60_command => cmd_R60_ne102, R62_command => cmd_R62_ne102, state => state_ne102, locking => ne102_locking);
	node_ne103 : node_44 port map(clock => clock, ocupation => ocupation(44), reset => reset, R21_command => cmd_R21_ne103, R28_command => cmd_R28_ne103, R30_command => cmd_R30_ne103, R46_command => cmd_R46_ne103, state => state_ne103, locking => ne103_locking);
	node_ne105 : node_45 port map(clock => clock, ocupation => ocupation(45), reset => reset, R9_command => cmd_R9_ne105, R19_command => cmd_R19_ne105, state => state_ne105, locking => ne105_locking);
	node_ne106 : node_46 port map(clock => clock, ocupation => ocupation(46), reset => reset, R10_command => cmd_R10_ne106, R22_command => cmd_R22_ne106, R32_command => cmd_R32_ne106, state => state_ne106, locking => ne106_locking);
	node_ne85 : node_47 port map(clock => clock, ocupation => ocupation(47), reset => reset, R6_command => cmd_R6_ne85, R78_command => cmd_R78_ne85, R79_command => cmd_R79_ne85, R80_command => cmd_R80_ne85, R86_command => cmd_R86_ne85, state => state_ne85, locking => ne85_locking);
	node_ne77 : node_48 port map(clock => clock, ocupation => ocupation(48), reset => reset, R65_command => cmd_R65_ne77, R81_command => cmd_R81_ne77, R82_command => cmd_R82_ne77, R89_command => cmd_R89_ne77, R90_command => cmd_R90_ne77, R91_command => cmd_R91_ne77, state => state_ne77, locking => ne77_locking);
	node_ne104 : node_49 port map(clock => clock, ocupation => ocupation(49), reset => reset, R14_command => cmd_R14_ne104, R87_command => cmd_R87_ne104, R88_command => cmd_R88_ne104, state => state_ne104, locking => ne104_locking);
	node_ne52 : node_50 port map(clock => clock, ocupation => ocupation(50), reset => reset, R3_command => cmd_R3_ne52, R42_command => cmd_R42_ne52, R44_command => cmd_R44_ne52, R45_command => cmd_R45_ne52, R81_command => cmd_R81_ne52, R91_command => cmd_R91_ne52, state => state_ne52, locking => ne52_locking);
	node_ne21 : node_51 port map(clock => clock, ocupation => ocupation(51), reset => reset, R14_command => cmd_R14_ne21, R35_command => cmd_R35_ne21, R36_command => cmd_R36_ne21, R37_command => cmd_R37_ne21, R66_command => cmd_R66_ne21, R83_command => cmd_R83_ne21, R88_command => cmd_R88_ne21, state => state_ne21, locking => ne21_locking);
	node_ne110 : node_52 port map(clock => clock, ocupation => ocupation(52), reset => reset, R54_command => cmd_R54_ne110, R56_command => cmd_R56_ne110, R58_command => cmd_R58_ne110, R59_command => cmd_R59_ne110, R84_command => cmd_R84_ne110, R85_command => cmd_R85_ne110, state => state_ne110, locking => ne110_locking);
	route_R1 : route_0 port map(clock => clock, routeRequest => routes_i(0), reset => reset, ne1_command => cmd_R1_ne1, ne1_state => state_ne1, ne1_lock => ne1_locking, T02_state => state_T02, T02_lock => T02_locking, T02_command => cmd_R1_T02, C78_state => state_C78, routeState => routes_o(0));
	route_R2 : route_1 port map(clock => clock, routeRequest => routes_i(1), reset => reset, ne7_command => cmd_R2_ne7, ne7_state => state_ne7, ne7_lock => ne7_locking, T06_state => state_T06, T06_lock => T06_locking, T06_command => cmd_R2_T06, J43_state => state_J43, routeState => routes_o(1));
	route_R3 : route_2 port map(clock => clock, routeRequest => routes_i(2), reset => reset, ne14_command => cmd_R3_ne14, ne14_state => state_ne14, ne14_lock => ne14_locking, ne52_command => cmd_R3_ne52, ne52_state => state_ne52, ne52_lock => ne52_locking, s69W04_command => cmd_R3_69W04, s69W04_state => state_69W04, s69W04_lock => s69W04_locking, T08_state => state_T08, T08_lock => T08_locking, T08_command => cmd_R3_T08, S146_state => state_S146, routeState => routes_o(2));
	route_R4 : route_3 port map(clock => clock, routeRequest => routes_i(3), reset => reset, ne47_command => cmd_R4_ne47, ne47_state => state_ne47, ne47_lock => ne47_locking, ne48_command => cmd_R4_ne48, ne48_state => state_ne48, ne48_lock => ne48_locking, s71W02_command => cmd_R4_71W02, s71W02_state => state_71W02, s71W02_lock => s71W02_locking, T12_state => state_T12, T12_lock => T12_locking, T12_command => cmd_R4_T12, L29_state => state_L29, routeState => routes_o(3));
	route_R5 : route_4 port map(clock => clock, routeRequest => routes_i(4), reset => reset, ne32_command => cmd_R5_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne82_command => cmd_R5_ne82, ne82_state => state_ne82, ne82_lock => ne82_locking, ne84_command => cmd_R5_ne84, ne84_state => state_ne84, ne84_lock => ne84_locking, Sw04_command => cmd_R5_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, Sw05_command => cmd_R5_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, T14_state => state_T14, T14_lock => T14_locking, T14_command => cmd_R5_T14, C100_state => state_C100, routeState => routes_o(4));
	route_R6 : route_5 port map(clock => clock, routeRequest => routes_i(5), reset => reset, ne44_command => cmd_R6_ne44, ne44_state => state_ne44, ne44_lock => ne44_locking, ne84_command => cmd_R6_ne84, ne84_state => state_ne84, ne84_lock => ne84_locking, ne100_command => cmd_R6_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne101_command => cmd_R6_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, ne85_command => cmd_R6_ne85, ne85_state => state_ne85, ne85_lock => ne85_locking, Sw05_command => cmd_R6_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, Sw41_command => cmd_R6_Sw41, Sw41_state => state_Sw41, Sw41_lock => Sw41_locking, T14_state => state_T14, T14_lock => T14_locking, T14_command => cmd_R6_T14, S105_state => state_S105, routeState => routes_o(5));
	route_R7 : route_6 port map(clock => clock, routeRequest => routes_i(6), reset => reset, ne30_command => cmd_R7_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne89_command => cmd_R7_ne89, ne89_state => state_ne89, ne89_lock => ne89_locking, Sw12_command => cmd_R7_Sw12, Sw12_state => state_Sw12, Sw12_lock => Sw12_locking, T20_state => state_T20, T20_lock => T20_locking, T20_command => cmd_R7_T20, S97_state => state_S97, routeState => routes_o(6));
	route_R8 : route_7 port map(clock => clock, routeRequest => routes_i(7), reset => reset, ne30_command => cmd_R8_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne90_command => cmd_R8_ne90, ne90_state => state_ne90, ne90_lock => ne90_locking, ne91_command => cmd_R8_ne91, ne91_state => state_ne91, ne91_lock => ne91_locking, Sw12_command => cmd_R8_Sw12, Sw12_state => state_Sw12, Sw12_lock => Sw12_locking, Sw13_command => cmd_R8_Sw13, Sw13_state => state_Sw13, Sw13_lock => Sw13_locking, T22_state => state_T22, T22_lock => T22_locking, T22_command => cmd_R8_T22, S97_state => state_S97, routeState => routes_o(7));
	route_R9 : route_8 port map(clock => clock, routeRequest => routes_i(8), reset => reset, ne96_command => cmd_R9_ne96, ne96_state => state_ne96, ne96_lock => ne96_locking, ne98_command => cmd_R9_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne105_command => cmd_R9_ne105, ne105_state => state_ne105, ne105_lock => ne105_locking, T24_state => state_T24, T24_lock => T24_locking, T24_command => cmd_R9_T24, P70_state => state_P70, routeState => routes_o(8));
	route_R10 : route_9 port map(clock => clock, routeRequest => routes_i(9), reset => reset, ne4_command => cmd_R10_ne4, ne4_state => state_ne4, ne4_lock => ne4_locking, ne106_command => cmd_R10_ne106, ne106_state => state_ne106, ne106_lock => ne106_locking, L25_state => state_L25, L25_lock => L25_locking, L25_command => cmd_R10_L25, L42_state => state_L42, routeState => routes_o(9));
	route_R11 : route_10 port map(clock => clock, routeRequest => routes_i(10), reset => reset, ne26_command => cmd_R11_ne26, ne26_state => state_ne26, ne26_lock => ne26_locking, ne65_command => cmd_R11_ne65, ne65_state => state_ne65, ne65_lock => ne65_locking, L27_state => state_L27, L27_lock => L27_locking, L27_command => cmd_R11_L27, L30_state => state_L30, routeState => routes_o(10));
	route_R12 : route_11 port map(clock => clock, routeRequest => routes_i(11), reset => reset, ne44_command => cmd_R12_ne44, ne44_state => state_ne44, ne44_lock => ne44_locking, ne101_command => cmd_R12_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, L28_state => state_L28, L28_lock => L28_locking, L28_command => cmd_R12_L28, L40_state => state_L40, routeState => routes_o(11));
	route_R13 : route_12 port map(clock => clock, routeRequest => routes_i(12), reset => reset, ne65_command => cmd_R13_ne65, ne65_state => state_ne65, ne65_lock => ne65_locking, ne102_command => cmd_R13_ne102, ne102_state => state_ne102, ne102_lock => ne102_locking, L30_state => state_L30, L30_lock => L30_locking, L30_command => cmd_R13_L30, C104_state => state_C104, routeState => routes_o(12));
	route_R14 : route_13 port map(clock => clock, routeRequest => routes_i(13), reset => reset, ne70_command => cmd_R14_ne70, ne70_state => state_ne70, ne70_lock => ne70_locking, ne104_command => cmd_R14_ne104, ne104_state => state_ne104, ne104_lock => ne104_locking, ne21_command => cmd_R14_ne21, ne21_state => state_ne21, ne21_lock => ne21_locking, Sw03_command => cmd_R14_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, L32_state => state_L32, L32_lock => L32_locking, L32_command => cmd_R14_L32, P73_state => state_P73, routeState => routes_o(13));
	route_R15 : route_14 port map(clock => clock, routeRequest => routes_i(14), reset => reset, ne78_command => cmd_R15_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, ne93_command => cmd_R15_ne93, ne93_state => state_ne93, ne93_lock => ne93_locking, L33_state => state_L33, L33_lock => L33_locking, L33_command => cmd_R15_L33, L34_state => state_L34, routeState => routes_o(14));
	route_R16 : route_15 port map(clock => clock, routeRequest => routes_i(15), reset => reset, ne93_command => cmd_R16_ne93, ne93_state => state_ne93, ne93_lock => ne93_locking, ne96_command => cmd_R16_ne96, ne96_state => state_ne96, ne96_lock => ne96_locking, L34_state => state_L34, L34_lock => L34_locking, L34_command => cmd_R16_L34, P71_state => state_P71, routeState => routes_o(15));
	route_R17 : route_16 port map(clock => clock, routeRequest => routes_i(16), reset => reset, ne95_command => cmd_R17_ne95, ne95_state => state_ne95, ne95_lock => ne95_locking, L35_state => state_L35, L35_lock => L35_locking, L35_command => cmd_R17_L35, X50_state => state_X50, routeState => routes_o(16));
	route_R18 : route_17 port map(clock => clock, routeRequest => routes_i(17), reset => reset, ne94_command => cmd_R18_ne94, ne94_state => state_ne94, ne94_lock => ne94_locking, ne97_command => cmd_R18_ne97, ne97_state => state_ne97, ne97_lock => ne97_locking, L37_state => state_L37, L37_lock => L37_locking, L37_command => cmd_R18_L37, S135_state => state_S135, routeState => routes_o(17));
	route_R19 : route_18 port map(clock => clock, routeRequest => routes_i(18), reset => reset, ne98_command => cmd_R19_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, ne105_command => cmd_R19_ne105, ne105_state => state_ne105, ne105_lock => ne105_locking, L38_state => state_L38, L38_lock => L38_locking, L38_command => cmd_R19_L38, T23_state => state_T23, routeState => routes_o(18));
	route_R20 : route_19 port map(clock => clock, routeRequest => routes_i(19), reset => reset, ne100_command => cmd_R20_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne101_command => cmd_R20_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, L40_state => state_L40, L40_lock => L40_locking, L40_command => cmd_R20_L40, S139_state => state_S139, routeState => routes_o(19));
	route_R21 : route_20 port map(clock => clock, routeRequest => routes_i(20), reset => reset, ne64_command => cmd_R21_ne64, ne64_state => state_ne64, ne64_lock => ne64_locking, ne103_command => cmd_R21_ne103, ne103_state => state_ne103, ne103_lock => ne103_locking, L41_state => state_L41, L41_lock => L41_locking, L41_command => cmd_R21_L41, S90_state => state_S90, routeState => routes_o(20));
	route_R22 : route_21 port map(clock => clock, routeRequest => routes_i(21), reset => reset, ne99_command => cmd_R22_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, ne106_command => cmd_R22_ne106, ne106_state => state_ne106, ne106_lock => ne106_locking, L42_state => state_L42, L42_lock => L42_locking, L42_command => cmd_R22_L42, P68_state => state_P68, routeState => routes_o(21));
	route_R23 : route_22 port map(clock => clock, routeRequest => routes_i(22), reset => reset, ne7_command => cmd_R23_ne7, ne7_state => state_ne7, ne7_lock => ne7_locking, ne9_command => cmd_R23_ne9, ne9_state => state_ne9, ne9_lock => ne9_locking, s68W02_command => cmd_R23_68W02, s68W02_state => state_68W02, s68W02_lock => s68W02_locking, J43_state => state_J43, J43_lock => J43_locking, J43_command => cmd_R23_J43, J46_state => state_J46, routeState => routes_o(22));
	route_R24 : route_23 port map(clock => clock, routeRequest => routes_i(23), reset => reset, ne9_command => cmd_R24_ne9, ne9_state => state_ne9, ne9_lock => ne9_locking, ne95_command => cmd_R24_ne95, ne95_state => state_ne95, ne95_lock => ne95_locking, J46_state => state_J46, J46_lock => J46_locking, J46_command => cmd_R24_J46, L35_state => state_L35, routeState => routes_o(23));
	route_R25 : route_24 port map(clock => clock, routeRequest => routes_i(24), reset => reset, ne59_command => cmd_R25_ne59, ne59_state => state_ne59, ne59_lock => ne59_locking, ne95_command => cmd_R25_ne95, ne95_state => state_ne95, ne95_lock => ne95_locking, Lc01_command => cmd_R25_Lc01, Lc01_state => state_Lc01, Lc01_lock => Lc01_locking, X50_state => state_X50, X50_lock => X50_locking, X50_command => cmd_R25_X50, S83_state => state_S83, routeState => routes_o(24));
	route_R26 : route_25 port map(clock => clock, routeRequest => routes_i(25), reset => reset, ne9_command => cmd_R26_ne9, ne9_state => state_ne9, ne9_lock => ne9_locking, ne95_command => cmd_R26_ne95, ne95_state => state_ne95, ne95_lock => ne95_locking, Lc01_command => cmd_R26_Lc01, Lc01_state => state_Lc01, Lc01_lock => Lc01_locking, X51_state => state_X51, X51_lock => X51_locking, X51_command => cmd_R26_X51, S80_state => state_S80, routeState => routes_o(25));
	route_R27 : route_26 port map(clock => clock, routeRequest => routes_i(26), reset => reset, ne23_command => cmd_R27_ne23, ne23_state => state_ne23, ne23_lock => ne23_locking, ne26_command => cmd_R27_ne26, ne26_state => state_ne26, ne26_lock => ne26_locking, s70W02_command => cmd_R27_70W02, s70W02_state => state_70W02, s70W02_lock => s70W02_locking, P60_state => state_P60, P60_lock => P60_locking, P60_command => cmd_R27_P60, L27_state => state_L27, routeState => routes_o(26));
	route_R28 : route_27 port map(clock => clock, routeRequest => routes_i(27), reset => reset, ne24_command => cmd_R28_ne24, ne24_state => state_ne24, ne24_lock => ne24_locking, ne64_command => cmd_R28_ne64, ne64_state => state_ne64, ne64_lock => ne64_locking, ne67_command => cmd_R28_ne67, ne67_state => state_ne67, ne67_lock => ne67_locking, ne103_command => cmd_R28_ne103, ne103_state => state_ne103, ne103_lock => ne103_locking, P63_state => state_P63, P63_lock => P63_locking, P63_command => cmd_R28_P63, P64_state => state_P64, routeState => routes_o(27));
	route_R29 : route_28 port map(clock => clock, routeRequest => routes_i(28), reset => reset, ne67_command => cmd_R29_ne67, ne67_state => state_ne67, ne67_lock => ne67_locking, ne70_command => cmd_R29_ne70, ne70_state => state_ne70, ne70_lock => ne70_locking, P64_state => state_P64, P64_lock => P64_locking, P64_command => cmd_R29_P64, L32_state => state_L32, routeState => routes_o(28));
	route_R30 : route_29 port map(clock => clock, routeRequest => routes_i(29), reset => reset, ne67_command => cmd_R30_ne67, ne67_state => state_ne67, ne67_lock => ne67_locking, ne103_command => cmd_R30_ne103, ne103_state => state_ne103, ne103_lock => ne103_locking, P65_state => state_P65, P65_lock => P65_locking, P65_command => cmd_R30_P65, L41_state => state_L41, routeState => routes_o(29));
	route_R31 : route_30 port map(clock => clock, routeRequest => routes_i(30), reset => reset, ne97_command => cmd_R31_ne97, ne97_state => state_ne97, ne97_lock => ne97_locking, ne99_command => cmd_R31_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, P68_state => state_P68, P68_lock => P68_locking, P68_command => cmd_R31_P68, L37_state => state_L37, routeState => routes_o(30));
	route_R32 : route_31 port map(clock => clock, routeRequest => routes_i(31), reset => reset, ne4_command => cmd_R32_ne4, ne4_state => state_ne4, ne4_lock => ne4_locking, ne99_command => cmd_R32_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, ne106_command => cmd_R32_ne106, ne106_state => state_ne106, ne106_lock => ne106_locking, P69_state => state_P69, P69_lock => P69_locking, P69_command => cmd_R32_P69, T03_state => state_T03, routeState => routes_o(31));
	route_R33 : route_32 port map(clock => clock, routeRequest => routes_i(32), reset => reset, ne78_command => cmd_R33_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, ne93_command => cmd_R33_ne93, ne93_state => state_ne93, ne93_lock => ne93_locking, ne96_command => cmd_R33_ne96, ne96_state => state_ne96, ne96_lock => ne96_locking, P70_state => state_P70, P70_lock => P70_locking, P70_command => cmd_R33_P70, S110_state => state_S110, routeState => routes_o(32));
	route_R34 : route_33 port map(clock => clock, routeRequest => routes_i(33), reset => reset, ne96_command => cmd_R34_ne96, ne96_state => state_ne96, ne96_lock => ne96_locking, ne98_command => cmd_R34_ne98, ne98_state => state_ne98, ne98_lock => ne98_locking, P71_state => state_P71, P71_lock => P71_locking, P71_command => cmd_R34_P71, L38_state => state_L38, routeState => routes_o(33));
	route_R35 : route_34 port map(clock => clock, routeRequest => routes_i(34), reset => reset, ne21_command => cmd_R35_ne21, ne21_state => state_ne21, ne21_lock => ne21_locking, P72_state => state_P72, P72_lock => P72_locking, P72_command => cmd_R35_P72, S144_state => state_S144, routeState => routes_o(34));
	route_R36 : route_35 port map(clock => clock, routeRequest => routes_i(35), reset => reset, ne78_command => cmd_R36_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, ne79_command => cmd_R36_ne79, ne79_state => state_ne79, ne79_lock => ne79_locking, ne21_command => cmd_R36_ne21, ne21_state => state_ne21, ne21_lock => ne21_locking, Sw06_command => cmd_R36_Sw06, Sw06_state => state_Sw06, Sw06_lock => Sw06_locking, Sw07_command => cmd_R36_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, P73_state => state_P73, P73_lock => P73_locking, P73_command => cmd_R36_P73, L33_state => state_L33, routeState => routes_o(35));
	route_R37 : route_36 port map(clock => clock, routeRequest => routes_i(36), reset => reset, ne94_command => cmd_R37_ne94, ne94_state => state_ne94, ne94_lock => ne94_locking, ne97_command => cmd_R37_ne97, ne97_state => state_ne97, ne97_lock => ne97_locking, ne99_command => cmd_R37_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, ne21_command => cmd_R37_ne21, ne21_state => state_ne21, ne21_lock => ne21_locking, Sw07_command => cmd_R37_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, P73_state => state_P73, P73_lock => P73_locking, P73_command => cmd_R37_P73, P69_state => state_P69, routeState => routes_o(36));
	route_R38 : route_37 port map(clock => clock, routeRequest => routes_i(37), reset => reset, ne1_command => cmd_R38_ne1, ne1_state => state_ne1, ne1_lock => ne1_locking, ne9_command => cmd_R38_ne9, ne9_state => state_ne9, ne9_lock => ne9_locking, s68W02_command => cmd_R38_68W02, s68W02_state => state_68W02, s68W02_lock => s68W02_locking, C78_state => state_C78, C78_lock => C78_locking, C78_command => cmd_R38_C78, J46_state => state_J46, routeState => routes_o(37));
	route_R39 : route_38 port map(clock => clock, routeRequest => routes_i(38), reset => reset, ne1_command => cmd_R39_ne1, ne1_state => state_ne1, ne1_lock => ne1_locking, ne9_command => cmd_R39_ne9, ne9_state => state_ne9, ne9_lock => ne9_locking, s68W02_command => cmd_R39_68W02, s68W02_state => state_68W02, s68W02_lock => s68W02_locking, S80_state => state_S80, S80_lock => S80_locking, S80_command => cmd_R39_S80, T01_state => state_T01, routeState => routes_o(38));
	route_R40 : route_39 port map(clock => clock, routeRequest => routes_i(39), reset => reset, ne7_command => cmd_R40_ne7, ne7_state => state_ne7, ne7_lock => ne7_locking, ne9_command => cmd_R40_ne9, ne9_state => state_ne9, ne9_lock => ne9_locking, s68W02_command => cmd_R40_68W02, s68W02_state => state_68W02, s68W02_lock => s68W02_locking, S80_state => state_S80, S80_lock => S80_locking, S80_command => cmd_R40_S80, T05_state => state_T05, routeState => routes_o(39));
	route_R41 : route_40 port map(clock => clock, routeRequest => routes_i(40), reset => reset, ne17_command => cmd_R41_ne17, ne17_state => state_ne17, ne17_lock => ne17_locking, ne59_command => cmd_R41_ne59, ne59_state => state_ne59, ne59_lock => ne59_locking, ne95_command => cmd_R41_ne95, ne95_state => state_ne95, ne95_lock => ne95_locking, s69W03_command => cmd_R41_69W03, s69W03_state => state_69W03, s69W03_lock => s69W03_locking, C82_state => state_C82, C82_lock => C82_locking, C82_command => cmd_R41_C82, X51_state => state_X51, routeState => routes_o(40));
	route_R42 : route_41 port map(clock => clock, routeRequest => routes_i(41), reset => reset, ne11_command => cmd_R42_ne11, ne11_state => state_ne11, ne11_lock => ne11_locking, ne59_command => cmd_R42_ne59, ne59_state => state_ne59, ne59_lock => ne59_locking, ne52_command => cmd_R42_ne52, ne52_state => state_ne52, ne52_lock => ne52_locking, s69W03_command => cmd_R42_69W03, s69W03_state => state_69W03, s69W03_lock => s69W03_locking, s69W04_command => cmd_R42_69W04, s69W04_state => state_69W04, s69W04_lock => s69W04_locking, S83_state => state_S83, S83_lock => S83_locking, S83_command => cmd_R42_S83, S146_state => state_S146, routeState => routes_o(41));
	route_R43 : route_42 port map(clock => clock, routeRequest => routes_i(42), reset => reset, ne17_command => cmd_R43_ne17, ne17_state => state_ne17, ne17_lock => ne17_locking, ne59_command => cmd_R43_ne59, ne59_state => state_ne59, ne59_lock => ne59_locking, s69W03_command => cmd_R43_69W03, s69W03_state => state_69W03, s69W03_lock => s69W03_locking, S83_state => state_S83, S83_lock => S83_locking, S83_command => cmd_R43_S83, C109_state => state_C109, routeState => routes_o(42));
	route_R44 : route_43 port map(clock => clock, routeRequest => routes_i(43), reset => reset, ne11_command => cmd_R44_ne11, ne11_state => state_ne11, ne11_lock => ne11_locking, ne59_command => cmd_R44_ne59, ne59_state => state_ne59, ne59_lock => ne59_locking, ne95_command => cmd_R44_ne95, ne95_state => state_ne95, ne95_lock => ne95_locking, ne52_command => cmd_R44_ne52, ne52_state => state_ne52, ne52_lock => ne52_locking, s69W03_command => cmd_R44_69W03, s69W03_state => state_69W03, s69W03_lock => s69W03_locking, s69W04_command => cmd_R44_69W04, s69W04_state => state_69W04, s69W04_lock => s69W04_locking, S86_state => state_S86, S86_lock => S86_locking, S86_command => cmd_R44_S86, X51_state => state_X51, routeState => routes_o(43));
	route_R45 : route_44 port map(clock => clock, routeRequest => routes_i(44), reset => reset, ne14_command => cmd_R45_ne14, ne14_state => state_ne14, ne14_lock => ne14_locking, ne52_command => cmd_R45_ne52, ne52_state => state_ne52, ne52_lock => ne52_locking, s69W04_command => cmd_R45_69W04, s69W04_state => state_69W04, s69W04_lock => s69W04_locking, S86_state => state_S86, S86_lock => S86_locking, S86_command => cmd_R45_S86, T07_state => state_T07, routeState => routes_o(44));
	route_R46 : route_45 port map(clock => clock, routeRequest => routes_i(45), reset => reset, ne23_command => cmd_R46_ne23, ne23_state => state_ne23, ne23_lock => ne23_locking, ne64_command => cmd_R46_ne64, ne64_state => state_ne64, ne64_lock => ne64_locking, ne67_command => cmd_R46_ne67, ne67_state => state_ne67, ne67_lock => ne67_locking, ne103_command => cmd_R46_ne103, ne103_state => state_ne103, ne103_lock => ne103_locking, B89_state => state_B89, B89_lock => B89_locking, B89_command => cmd_R46_B89, P64_state => state_P64, routeState => routes_o(45));
	route_R47 : route_46 port map(clock => clock, routeRequest => routes_i(46), reset => reset, ne23_command => cmd_R47_ne23, ne23_state => state_ne23, ne23_lock => ne23_locking, ne64_command => cmd_R47_ne64, ne64_state => state_ne64, ne64_lock => ne64_locking, s70W01_command => cmd_R47_70W01, s70W01_state => state_70W01, s70W01_lock => s70W01_locking, S90_state => state_S90, S90_lock => S90_locking, S90_command => cmd_R47_S90, P60_state => state_P60, routeState => routes_o(46));
	route_R48 : route_47 port map(clock => clock, routeRequest => routes_i(47), reset => reset, ne24_command => cmd_R48_ne24, ne24_state => state_ne24, ne24_lock => ne24_locking, ne64_command => cmd_R48_ne64, ne64_state => state_ne64, ne64_lock => ne64_locking, s70W01_command => cmd_R48_70W01, s70W01_state => state_70W01, s70W01_lock => s70W01_locking, S90_state => state_S90, S90_lock => S90_locking, S90_command => cmd_R48_S90, B92_state => state_B92, routeState => routes_o(47));
	route_R49 : route_48 port map(clock => clock, routeRequest => routes_i(48), reset => reset, ne24_command => cmd_R49_ne24, ne24_state => state_ne24, ne24_lock => ne24_locking, ne26_command => cmd_R49_ne26, ne26_state => state_ne26, ne26_lock => ne26_locking, s70W02_command => cmd_R49_70W02, s70W02_state => state_70W02, s70W02_lock => s70W02_locking, B92_state => state_B92, B92_lock => B92_locking, B92_command => cmd_R49_B92, L27_state => state_L27, routeState => routes_o(48));
	route_R50 : route_49 port map(clock => clock, routeRequest => routes_i(49), reset => reset, ne23_command => cmd_R50_ne23, ne23_state => state_ne23, ne23_lock => ne23_locking, ne26_command => cmd_R50_ne26, ne26_state => state_ne26, ne26_lock => ne26_locking, s70W02_command => cmd_R50_70W02, s70W02_state => state_70W02, s70W02_lock => s70W02_locking, S93_state => state_S93, S93_lock => S93_locking, S93_command => cmd_R50_S93, B89_state => state_B89, routeState => routes_o(49));
	route_R51 : route_50 port map(clock => clock, routeRequest => routes_i(50), reset => reset, ne24_command => cmd_R51_ne24, ne24_state => state_ne24, ne24_lock => ne24_locking, ne26_command => cmd_R51_ne26, ne26_state => state_ne26, ne26_lock => ne26_locking, s70W02_command => cmd_R51_70W02, s70W02_state => state_70W02, s70W02_lock => s70W02_locking, S93_state => state_S93, S93_lock => S93_locking, S93_command => cmd_R51_S93, P63_state => state_P63, routeState => routes_o(50));
	route_R52 : route_51 port map(clock => clock, routeRequest => routes_i(51), reset => reset, ne30_command => cmd_R52_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne83_command => cmd_R52_ne83, ne83_state => state_ne83, ne83_lock => ne83_locking, Sw08_command => cmd_R52_Sw08, Sw08_state => state_Sw08, Sw08_lock => Sw08_locking, C95_state => state_C95, C95_lock => C95_locking, C95_command => cmd_R52_C95, S122_state => state_S122, routeState => routes_o(51));
	route_R53 : route_52 port map(clock => clock, routeRequest => routes_i(52), reset => reset, ne29_command => cmd_R53_ne29, ne29_state => state_ne29, ne29_lock => ne29_locking, ne30_command => cmd_R53_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, Sw08_command => cmd_R53_Sw08, Sw08_state => state_Sw08, Sw08_lock => Sw08_locking, B96_state => state_B96, B96_lock => B96_locking, B96_command => cmd_R53_B96, S122_state => state_S122, routeState => routes_o(52));
	route_R54 : route_53 port map(clock => clock, routeRequest => routes_i(53), reset => reset, ne29_command => cmd_R54_ne29, ne29_state => state_ne29, ne29_lock => ne29_locking, ne30_command => cmd_R54_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne110_command => cmd_R54_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, Sw08_command => cmd_R54_Sw08, Sw08_state => state_Sw08, Sw08_lock => Sw08_locking, Sw09_command => cmd_R54_Sw09, Sw09_state => state_Sw09, Sw09_lock => Sw09_locking, S97_state => state_S97, S97_lock => S97_locking, S97_command => cmd_R54_S97, C138_state => state_C138, routeState => routes_o(53));
	route_R55 : route_54 port map(clock => clock, routeRequest => routes_i(54), reset => reset, ne30_command => cmd_R55_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne83_command => cmd_R55_ne83, ne83_state => state_ne83, ne83_lock => ne83_locking, Sw08_command => cmd_R55_Sw08, Sw08_state => state_Sw08, Sw08_lock => Sw08_locking, S97_state => state_S97, S97_lock => S97_locking, S97_command => cmd_R55_S97, C114_state => state_C114, routeState => routes_o(54));
	route_R56 : route_55 port map(clock => clock, routeRequest => routes_i(55), reset => reset, ne32_command => cmd_R56_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne110_command => cmd_R56_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, Sw09_command => cmd_R56_Sw09, Sw09_state => state_Sw09, Sw09_lock => Sw09_locking, C100_state => state_C100, C100_lock => C100_locking, C100_command => cmd_R56_C100, C138_state => state_C138, routeState => routes_o(55));
	route_R57 : route_56 port map(clock => clock, routeRequest => routes_i(56), reset => reset, ne29_command => cmd_R57_ne29, ne29_state => state_ne29, ne29_lock => ne29_locking, B101_state => state_B101, B101_lock => B101_locking, B101_command => cmd_R57_B101, B96_state => state_B96, routeState => routes_o(56));
	route_R58 : route_57 port map(clock => clock, routeRequest => routes_i(57), reset => reset, ne32_command => cmd_R58_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne110_command => cmd_R58_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, Sw09_command => cmd_R58_Sw09, Sw09_state => state_Sw09, Sw09_lock => Sw09_locking, S102_state => state_S102, S102_lock => S102_locking, S102_command => cmd_R58_S102, S115_state => state_S115, routeState => routes_o(57));
	route_R59 : route_58 port map(clock => clock, routeRequest => routes_i(58), reset => reset, ne29_command => cmd_R59_ne29, ne29_state => state_ne29, ne29_lock => ne29_locking, ne110_command => cmd_R59_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, Sw09_command => cmd_R59_Sw09, Sw09_state => state_Sw09, Sw09_lock => Sw09_locking, S102_state => state_S102, S102_lock => S102_locking, S102_command => cmd_R59_S102, B101_state => state_B101, routeState => routes_o(58));
	route_R60 : route_59 port map(clock => clock, routeRequest => routes_i(59), reset => reset, ne44_command => cmd_R60_ne44, ne44_state => state_ne44, ne44_lock => ne44_locking, ne102_command => cmd_R60_ne102, ne102_state => state_ne102, ne102_lock => ne102_locking, s71W01_command => cmd_R60_71W01, s71W01_state => state_71W01, s71W01_lock => s71W01_locking, C104_state => state_C104, C104_lock => C104_locking, C104_command => cmd_R60_C104, L28_state => state_L28, routeState => routes_o(59));
	route_R61 : route_60 port map(clock => clock, routeRequest => routes_i(60), reset => reset, ne43_command => cmd_R61_ne43, ne43_state => state_ne43, ne43_lock => ne43_locking, ne44_command => cmd_R61_ne44, ne44_state => state_ne44, ne44_lock => ne44_locking, ne48_command => cmd_R61_ne48, ne48_state => state_ne48, ne48_lock => ne48_locking, s71W01_command => cmd_R61_71W01, s71W01_state => state_71W01, s71W01_lock => s71W01_locking, s71W02_command => cmd_R61_71W02, s71W02_state => state_71W02, s71W02_lock => s71W02_locking, S105_state => state_S105, S105_lock => S105_locking, S105_command => cmd_R61_S105, L29_state => state_L29, routeState => routes_o(60));
	route_R62 : route_61 port map(clock => clock, routeRequest => routes_i(61), reset => reset, ne26_command => cmd_R62_ne26, ne26_state => state_ne26, ne26_lock => ne26_locking, ne44_command => cmd_R62_ne44, ne44_state => state_ne44, ne44_lock => ne44_locking, ne65_command => cmd_R62_ne65, ne65_state => state_ne65, ne65_lock => ne65_locking, ne102_command => cmd_R62_ne102, ne102_state => state_ne102, ne102_lock => ne102_locking, s71W01_command => cmd_R62_71W01, s71W01_state => state_71W01, s71W01_lock => s71W01_locking, S105_state => state_S105, S105_lock => S105_locking, S105_command => cmd_R62_S105, S93_state => state_S93, routeState => routes_o(61));
	route_R63 : route_62 port map(clock => clock, routeRequest => routes_i(62), reset => reset, ne17_command => cmd_R63_ne17, ne17_state => state_ne17, ne17_lock => ne17_locking, ne78_command => cmd_R63_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, Sw06_command => cmd_R63_Sw06, Sw06_state => state_Sw06, Sw06_lock => Sw06_locking, C109_state => state_C109, C109_lock => C109_locking, C109_command => cmd_R63_C109, L33_state => state_L33, routeState => routes_o(62));
	route_R64 : route_63 port map(clock => clock, routeRequest => routes_i(63), reset => reset, ne17_command => cmd_R64_ne17, ne17_state => state_ne17, ne17_lock => ne17_locking, ne78_command => cmd_R64_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, Sw06_command => cmd_R64_Sw06, Sw06_state => state_Sw06, Sw06_lock => Sw06_locking, S110_state => state_S110, S110_lock => S110_locking, S110_command => cmd_R64_S110, C82_state => state_C82, routeState => routes_o(63));
	route_R65 : route_64 port map(clock => clock, routeRequest => routes_i(64), reset => reset, ne78_command => cmd_R65_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, ne79_command => cmd_R65_ne79, ne79_state => state_ne79, ne79_lock => ne79_locking, ne77_command => cmd_R65_ne77, ne77_state => state_ne77, ne77_lock => ne77_locking, Sw06_command => cmd_R65_Sw06, Sw06_state => state_Sw06, Sw06_lock => Sw06_locking, Sw07_command => cmd_R65_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, S110_state => state_S110, S110_lock => S110_locking, S110_command => cmd_R65_S110, B133_state => state_B133, routeState => routes_o(64));
	route_R66 : route_65 port map(clock => clock, routeRequest => routes_i(65), reset => reset, ne78_command => cmd_R66_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, ne79_command => cmd_R66_ne79, ne79_state => state_ne79, ne79_lock => ne79_locking, ne21_command => cmd_R66_ne21, ne21_state => state_ne21, ne21_lock => ne21_locking, Sw06_command => cmd_R66_Sw06, Sw06_state => state_Sw06, Sw06_lock => Sw06_locking, Sw07_command => cmd_R66_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, S110_state => state_S110, S110_lock => S110_locking, S110_command => cmd_R66_S110, P72_state => state_P72, routeState => routes_o(65));
	route_R67 : route_66 port map(clock => clock, routeRequest => routes_i(66), reset => reset, ne32_command => cmd_R67_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne83_command => cmd_R67_ne83, ne83_state => state_ne83, ne83_lock => ne83_locking, Sw04_command => cmd_R67_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, C114_state => state_C114, C114_lock => C114_locking, C114_command => cmd_R67_C114, C100_state => state_C100, routeState => routes_o(66));
	route_R68 : route_67 port map(clock => clock, routeRequest => routes_i(67), reset => reset, ne32_command => cmd_R68_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne83_command => cmd_R68_ne83, ne83_state => state_ne83, ne83_lock => ne83_locking, Sw04_command => cmd_R68_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, S115_state => state_S115, S115_lock => S115_locking, S115_command => cmd_R68_S115, C95_state => state_C95, routeState => routes_o(67));
	route_R69 : route_68 port map(clock => clock, routeRequest => routes_i(68), reset => reset, ne32_command => cmd_R69_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne41_command => cmd_R69_ne41, ne41_state => state_ne41, ne41_lock => ne41_locking, ne82_command => cmd_R69_ne82, ne82_state => state_ne82, ne82_lock => ne82_locking, Sw04_command => cmd_R69_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, Sw05_command => cmd_R69_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, S115_state => state_S115, S115_lock => S115_locking, S115_command => cmd_R69_S115, P58_state => state_P58, routeState => routes_o(68));
	route_R70 : route_69 port map(clock => clock, routeRequest => routes_i(69), reset => reset, ne32_command => cmd_R70_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne82_command => cmd_R70_ne82, ne82_state => state_ne82, ne82_lock => ne82_locking, ne84_command => cmd_R70_ne84, ne84_state => state_ne84, ne84_lock => ne84_locking, Sw04_command => cmd_R70_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, Sw05_command => cmd_R70_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, S115_state => state_S115, S115_lock => S115_locking, S115_command => cmd_R70_S115, T13_state => state_T13, routeState => routes_o(69));
	route_R71 : route_70 port map(clock => clock, routeRequest => routes_i(70), reset => reset, ne86_command => cmd_R71_ne86, ne86_state => state_ne86, ne86_lock => ne86_locking, ne88_command => cmd_R71_ne88, ne88_state => state_ne88, ne88_lock => ne88_locking, Sw11_command => cmd_R71_Sw11, Sw11_state => state_Sw11, Sw11_lock => Sw11_locking, C118_state => state_C118, C118_lock => C118_locking, C118_command => cmd_R71_C118, T15_state => state_T15, routeState => routes_o(70));
	route_R72 : route_71 port map(clock => clock, routeRequest => routes_i(71), reset => reset, ne86_command => cmd_R72_ne86, ne86_state => state_ne86, ne86_lock => ne86_locking, ne88_command => cmd_R72_ne88, ne88_state => state_ne88, ne88_lock => ne88_locking, Sw11_command => cmd_R72_Sw11, Sw11_state => state_Sw11, Sw11_lock => Sw11_locking, S119_state => state_S119, S119_lock => S119_locking, S119_command => cmd_R72_S119, T17_state => state_T17, routeState => routes_o(71));
	route_R73 : route_72 port map(clock => clock, routeRequest => routes_i(72), reset => reset, ne30_command => cmd_R73_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne86_command => cmd_R73_ne86, ne86_state => state_ne86, ne86_lock => ne86_locking, ne87_command => cmd_R73_ne87, ne87_state => state_ne87, ne87_lock => ne87_locking, ne91_command => cmd_R73_ne91, ne91_state => state_ne91, ne91_lock => ne91_locking, Sw11_command => cmd_R73_Sw11, Sw11_state => state_Sw11, Sw11_lock => Sw11_locking, Sw12_command => cmd_R73_Sw12, Sw12_state => state_Sw12, Sw12_lock => Sw12_locking, Sw13_command => cmd_R73_Sw13, Sw13_state => state_Sw13, Sw13_lock => Sw13_locking, S119_state => state_S119, S119_lock => S119_locking, S119_command => cmd_R73_S119, S97_state => state_S97, routeState => routes_o(72));
	route_R74 : route_73 port map(clock => clock, routeRequest => routes_i(73), reset => reset, ne30_command => cmd_R74_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne89_command => cmd_R74_ne89, ne89_state => state_ne89, ne89_lock => ne89_locking, Sw12_command => cmd_R74_Sw12, Sw12_state => state_Sw12, Sw12_lock => Sw12_locking, S122_state => state_S122, S122_lock => S122_locking, S122_command => cmd_R74_S122, T19_state => state_T19, routeState => routes_o(73));
	route_R75 : route_74 port map(clock => clock, routeRequest => routes_i(74), reset => reset, ne30_command => cmd_R75_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne86_command => cmd_R75_ne86, ne86_state => state_ne86, ne86_lock => ne86_locking, ne87_command => cmd_R75_ne87, ne87_state => state_ne87, ne87_lock => ne87_locking, ne91_command => cmd_R75_ne91, ne91_state => state_ne91, ne91_lock => ne91_locking, Sw11_command => cmd_R75_Sw11, Sw11_state => state_Sw11, Sw11_lock => Sw11_locking, Sw12_command => cmd_R75_Sw12, Sw12_state => state_Sw12, Sw12_lock => Sw12_locking, Sw13_command => cmd_R75_Sw13, Sw13_state => state_Sw13, Sw13_lock => Sw13_locking, S122_state => state_S122, S122_lock => S122_locking, S122_command => cmd_R75_S122, T15_state => state_T15, routeState => routes_o(74));
	route_R76 : route_75 port map(clock => clock, routeRequest => routes_i(75), reset => reset, ne30_command => cmd_R76_ne30, ne30_state => state_ne30, ne30_lock => ne30_locking, ne90_command => cmd_R76_ne90, ne90_state => state_ne90, ne90_lock => ne90_locking, ne91_command => cmd_R76_ne91, ne91_state => state_ne91, ne91_lock => ne91_locking, Sw12_command => cmd_R76_Sw12, Sw12_state => state_Sw12, Sw12_lock => Sw12_locking, Sw13_command => cmd_R76_Sw13, Sw13_state => state_Sw13, Sw13_lock => Sw13_locking, S122_state => state_S122, S122_lock => S122_locking, S122_command => cmd_R76_S122, T21_state => state_T21, routeState => routes_o(75));
	route_R77 : route_76 port map(clock => clock, routeRequest => routes_i(76), reset => reset, ne32_command => cmd_R77_ne32, ne32_state => state_ne32, ne32_lock => ne32_locking, ne41_command => cmd_R77_ne41, ne41_state => state_ne41, ne41_lock => ne41_locking, ne82_command => cmd_R77_ne82, ne82_state => state_ne82, ne82_lock => ne82_locking, Sw04_command => cmd_R77_Sw04, Sw04_state => state_Sw04, Sw04_lock => Sw04_locking, Sw05_command => cmd_R77_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, B130_state => state_B130, B130_lock => B130_locking, B130_command => cmd_R77_B130, C100_state => state_C100, routeState => routes_o(76));
	route_R78 : route_77 port map(clock => clock, routeRequest => routes_i(77), reset => reset, ne41_command => cmd_R78_ne41, ne41_state => state_ne41, ne41_lock => ne41_locking, ne44_command => cmd_R78_ne44, ne44_state => state_ne44, ne44_lock => ne44_locking, ne100_command => cmd_R78_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne101_command => cmd_R78_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, ne85_command => cmd_R78_ne85, ne85_state => state_ne85, ne85_lock => ne85_locking, Sw05_command => cmd_R78_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, Sw41_command => cmd_R78_Sw41, Sw41_state => state_Sw41, Sw41_lock => Sw41_locking, B130_state => state_B130, B130_lock => B130_locking, B130_command => cmd_R78_B130, S105_state => state_S105, routeState => routes_o(77));
	route_R79 : route_78 port map(clock => clock, routeRequest => routes_i(78), reset => reset, ne41_command => cmd_R79_ne41, ne41_state => state_ne41, ne41_lock => ne41_locking, ne85_command => cmd_R79_ne85, ne85_state => state_ne85, ne85_lock => ne85_locking, Sw05_command => cmd_R79_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, S131_state => state_S131, S131_lock => S131_locking, S131_command => cmd_R79_S131, P58_state => state_P58, routeState => routes_o(78));
	route_R80 : route_79 port map(clock => clock, routeRequest => routes_i(79), reset => reset, ne84_command => cmd_R80_ne84, ne84_state => state_ne84, ne84_lock => ne84_locking, ne85_command => cmd_R80_ne85, ne85_state => state_ne85, ne85_lock => ne85_locking, Sw05_command => cmd_R80_Sw05, Sw05_state => state_Sw05, Sw05_lock => Sw05_locking, S131_state => state_S131, S131_lock => S131_locking, S131_command => cmd_R80_S131, T13_state => state_T13, routeState => routes_o(79));
	route_R81 : route_80 port map(clock => clock, routeRequest => routes_i(80), reset => reset, ne77_command => cmd_R81_ne77, ne77_state => state_ne77, ne77_lock => ne77_locking, ne52_command => cmd_R81_ne52, ne52_state => state_ne52, ne52_lock => ne52_locking, Sw03_command => cmd_R81_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, B133_state => state_B133, B133_lock => B133_locking, B133_command => cmd_R81_B133, S86_state => state_S86, routeState => routes_o(80));
	route_R82 : route_81 port map(clock => clock, routeRequest => routes_i(81), reset => reset, ne94_command => cmd_R82_ne94, ne94_state => state_ne94, ne94_lock => ne94_locking, ne77_command => cmd_R82_ne77, ne77_state => state_ne77, ne77_lock => ne77_locking, Sw07_command => cmd_R82_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, S135_state => state_S135, S135_lock => S135_locking, S135_command => cmd_R82_S135, B133_state => state_B133, routeState => routes_o(81));
	route_R83 : route_82 port map(clock => clock, routeRequest => routes_i(82), reset => reset, ne94_command => cmd_R83_ne94, ne94_state => state_ne94, ne94_lock => ne94_locking, ne21_command => cmd_R83_ne21, ne21_state => state_ne21, ne21_lock => ne21_locking, Sw07_command => cmd_R83_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, S135_state => state_S135, S135_lock => S135_locking, S135_command => cmd_R83_S135, P72_state => state_P72, routeState => routes_o(82));
	route_R84 : route_83 port map(clock => clock, routeRequest => routes_i(83), reset => reset, ne44_command => cmd_R84_ne44, ne44_state => state_ne44, ne44_lock => ne44_locking, ne100_command => cmd_R84_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne101_command => cmd_R84_ne101, ne101_state => state_ne101, ne101_lock => ne101_locking, ne110_command => cmd_R84_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, Sw41_command => cmd_R84_Sw41, Sw41_state => state_Sw41, Sw41_lock => Sw41_locking, C138_state => state_C138, C138_lock => C138_locking, C138_command => cmd_R84_C138, S105_state => state_S105, routeState => routes_o(83));
	route_R85 : route_84 port map(clock => clock, routeRequest => routes_i(84), reset => reset, ne100_command => cmd_R85_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne110_command => cmd_R85_ne110, ne110_state => state_ne110, ne110_lock => ne110_locking, Sw41_command => cmd_R85_Sw41, Sw41_state => state_Sw41, Sw41_lock => Sw41_locking, S139_state => state_S139, S139_lock => S139_locking, S139_command => cmd_R85_S139, S102_state => state_S102, routeState => routes_o(84));
	route_R86 : route_85 port map(clock => clock, routeRequest => routes_i(85), reset => reset, ne100_command => cmd_R86_ne100, ne100_state => state_ne100, ne100_lock => ne100_locking, ne85_command => cmd_R86_ne85, ne85_state => state_ne85, ne85_lock => ne85_locking, Sw41_command => cmd_R86_Sw41, Sw41_state => state_Sw41, Sw41_lock => Sw41_locking, S139_state => state_S139, S139_lock => S139_locking, S139_command => cmd_R86_S139, S131_state => state_S131, routeState => routes_o(85));
	route_R87 : route_86 port map(clock => clock, routeRequest => routes_i(86), reset => reset, ne70_command => cmd_R87_ne70, ne70_state => state_ne70, ne70_lock => ne70_locking, ne104_command => cmd_R87_ne104, ne104_state => state_ne104, ne104_lock => ne104_locking, B143_state => state_B143, B143_lock => B143_locking, B143_command => cmd_R87_B143, L32_state => state_L32, routeState => routes_o(86));
	route_R88 : route_87 port map(clock => clock, routeRequest => routes_i(87), reset => reset, ne104_command => cmd_R88_ne104, ne104_state => state_ne104, ne104_lock => ne104_locking, ne21_command => cmd_R88_ne21, ne21_state => state_ne21, ne21_lock => ne21_locking, Sw03_command => cmd_R88_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, S144_state => state_S144, S144_lock => S144_locking, S144_command => cmd_R88_S144, B143_state => state_B143, routeState => routes_o(87));
	route_R89 : route_88 port map(clock => clock, routeRequest => routes_i(88), reset => reset, ne78_command => cmd_R89_ne78, ne78_state => state_ne78, ne78_lock => ne78_locking, ne79_command => cmd_R89_ne79, ne79_state => state_ne79, ne79_lock => ne79_locking, ne77_command => cmd_R89_ne77, ne77_state => state_ne77, ne77_lock => ne77_locking, Sw06_command => cmd_R89_Sw06, Sw06_state => state_Sw06, Sw06_lock => Sw06_locking, Sw07_command => cmd_R89_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, B145_state => state_B145, B145_lock => B145_locking, B145_command => cmd_R89_B145, L33_state => state_L33, routeState => routes_o(88));
	route_R90 : route_89 port map(clock => clock, routeRequest => routes_i(89), reset => reset, ne94_command => cmd_R90_ne94, ne94_state => state_ne94, ne94_lock => ne94_locking, ne97_command => cmd_R90_ne97, ne97_state => state_ne97, ne97_lock => ne97_locking, ne99_command => cmd_R90_ne99, ne99_state => state_ne99, ne99_lock => ne99_locking, ne77_command => cmd_R90_ne77, ne77_state => state_ne77, ne77_lock => ne77_locking, Sw07_command => cmd_R90_Sw07, Sw07_state => state_Sw07, Sw07_lock => Sw07_locking, B145_state => state_B145, B145_lock => B145_locking, B145_command => cmd_R90_B145, P69_state => state_P69, routeState => routes_o(89));
	route_R91 : route_90 port map(clock => clock, routeRequest => routes_i(90), reset => reset, ne77_command => cmd_R91_ne77, ne77_state => state_ne77, ne77_lock => ne77_locking, ne52_command => cmd_R91_ne52, ne52_state => state_ne52, ne52_lock => ne52_locking, Sw03_command => cmd_R91_Sw03, Sw03_state => state_Sw03, Sw03_lock => Sw03_locking, S146_state => state_S146, S146_lock => S146_locking, S146_command => cmd_R91_S146, B145_state => state_B145, routeState => routes_o(90));
	processed <= processing;
end Behavioral;