--  network.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
--Declare the package
use work.my_package.all;
	entity network is
		generic(
			N_TRACKCIRCUITS : natural := 53;
			N_ROUTES : natural := 91;
			N_SIGNALS : natural := 82;
			N_LEVELCROSSINGS : natural := 1;
			N_SINGLESWITCHES : natural := 15;
			N_DOUBLESWITCHES : natural := 2;
			N_SCISSORCROSSINGS : natural := 1;
			N : natural := 245
		);
		port(
			clock : in std_logic;
			processing : in std_logic;
			processed : out std_logic;
			tracks_i : in hex_array(N_TRACKCIRCUITS-1 downto 0);
			tracks_o : out hex_array(N_TRACKCIRCUITS-1 downto 0);
			signals_i : in hex_array(N_SIGNALS-1 downto 0);
			signals_o : out hex_array(N_SIGNALS-1 downto 0);
			routes_i : in hex_array(N_ROUTES-1 downto 0);
			routes_o : out hex_array(N_ROUTES-1 downto 0);
			levelCrossings_i : in hex_char;
			levelCrossings_o : out hex_char;
			singleSwitches_i : in hex_array(N_SINGLESWITCHES-1 downto 0);
			singleSwitches_o : out hex_array(N_SINGLESWITCHES-1 downto 0);
			scissorCrossings_i : in hex_char;
			scissorCrossings_o : out hex_char;
			doubleSwitches_i : in hex_array(N_DOUBLESWITCHES-1 downto 0);
			doubleSwitches_o : out hex_array(N_DOUBLESWITCHES-1 downto 0);
			reset : in std_logic
		);
	end entity network;
architecture Behavioral of network is
	component levelCrossing_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			track_ne95 : in hex_char;
			track_ne9 : in hex_char;
			track_ne59 : in hex_char;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			R41_command : in routeCommands;
			R44_command : in routeCommands;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component levelCrossing_0;
	component singleSwitch_0 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R23_command : in routeCommands := RELEASE;
			R38_command : in routeCommands := RELEASE;
			R39_command : in routeCommands := RELEASE;
			R40_command : in routeCommands := RELEASE;
			R1_command : in routeCommands := RELEASE;
			R2_command : in routeCommands := RELEASE;
			R26_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_0;
	component singleSwitch_1 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R41_command : in routeCommands := RELEASE;
			R42_command : in routeCommands := RELEASE;
			R43_command : in routeCommands := RELEASE;
			R44_command : in routeCommands := RELEASE;
			R64_command : in routeCommands := RELEASE;
			R25_command : in routeCommands := RELEASE;
			R81_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_1;
	component singleSwitch_2 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R3_command : in routeCommands := RELEASE;
			R42_command : in routeCommands := RELEASE;
			R44_command : in routeCommands := RELEASE;
			R45_command : in routeCommands := RELEASE;
			R25_command : in routeCommands := RELEASE;
			R81_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_2;
	component singleSwitch_3 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R36_command : in routeCommands := RELEASE;
			R63_command : in routeCommands := RELEASE;
			R64_command : in routeCommands := RELEASE;
			R65_command : in routeCommands := RELEASE;
			R66_command : in routeCommands := RELEASE;
			R89_command : in routeCommands := RELEASE;
			R43_command : in routeCommands := RELEASE;
			R14_command : in routeCommands := RELEASE;
			R33_command : in routeCommands := RELEASE;
			R91_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_3;
	component singleSwitch_4 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R47_command : in routeCommands := RELEASE;
			R48_command : in routeCommands := RELEASE;
			R21_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_4;
	component singleSwitch_5 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R27_command : in routeCommands := RELEASE;
			R49_command : in routeCommands := RELEASE;
			R50_command : in routeCommands := RELEASE;
			R51_command : in routeCommands := RELEASE;
			R62_command : in routeCommands := RELEASE;
			R47_command : in routeCommands := RELEASE;
			R48_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_5;
	component singleSwitch_6 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R52_command : in routeCommands := RELEASE;
			R53_command : in routeCommands := RELEASE;
			R54_command : in routeCommands := RELEASE;
			R55_command : in routeCommands := RELEASE;
			R57_command : in routeCommands := RELEASE;
			R68_command : in routeCommands := RELEASE;
			R73_command : in routeCommands := RELEASE;
			R7_command : in routeCommands := RELEASE;
			R8_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_6;
	component singleSwitch_7 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R54_command : in routeCommands := RELEASE;
			R56_command : in routeCommands := RELEASE;
			R58_command : in routeCommands := RELEASE;
			R59_command : in routeCommands := RELEASE;
			R77_command : in routeCommands := RELEASE;
			R67_command : in routeCommands := RELEASE;
			R5_command : in routeCommands := RELEASE;
			R73_command : in routeCommands := RELEASE;
			R7_command : in routeCommands := RELEASE;
			R8_command : in routeCommands := RELEASE;
			R85_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_7;
	component singleSwitch_8 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R7_command : in routeCommands := RELEASE;
			R8_command : in routeCommands := RELEASE;
			R73_command : in routeCommands := RELEASE;
			R74_command : in routeCommands := RELEASE;
			R75_command : in routeCommands := RELEASE;
			R76_command : in routeCommands := RELEASE;
			R53_command : in routeCommands := RELEASE;
			R52_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_8;
	component singleSwitch_9 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R5_command : in routeCommands := RELEASE;
			R67_command : in routeCommands := RELEASE;
			R68_command : in routeCommands := RELEASE;
			R69_command : in routeCommands := RELEASE;
			R70_command : in routeCommands := RELEASE;
			R77_command : in routeCommands := RELEASE;
			R55_command : in routeCommands := RELEASE;
			R58_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_9;
	component singleSwitch_10 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R60_command : in routeCommands := RELEASE;
			R61_command : in routeCommands := RELEASE;
			R62_command : in routeCommands := RELEASE;
			R78_command : in routeCommands := RELEASE;
			R13_command : in routeCommands := RELEASE;
			R6_command : in routeCommands := RELEASE;
			R84_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_10;
	component singleSwitch_11 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R4_command : in routeCommands := RELEASE;
			R61_command : in routeCommands := RELEASE;
			R78_command : in routeCommands := RELEASE;
			R6_command : in routeCommands := RELEASE;
			R84_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_11;
	component singleSwitch_12 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R71_command : in routeCommands := RELEASE;
			R72_command : in routeCommands := RELEASE;
			R73_command : in routeCommands := RELEASE;
			R75_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_12;
	component singleSwitch_13 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R8_command : in routeCommands := RELEASE;
			R73_command : in routeCommands := RELEASE;
			R75_command : in routeCommands := RELEASE;
			R76_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_13;
	component singleSwitch_14 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R6_command : in routeCommands := RELEASE;
			R78_command : in routeCommands := RELEASE;
			R84_command : in routeCommands := RELEASE;
			R85_command : in routeCommands := RELEASE;
			R86_command : in routeCommands := RELEASE;
			R54_command : in routeCommands := RELEASE;
			R56_command : in routeCommands := RELEASE;
			R20_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component singleSwitch_14;
	component scissorCrossing_0 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R14_command : in routeCommands := RELEASE;
			R81_command : in routeCommands := RELEASE;
			R88_command : in routeCommands := RELEASE;
			R91_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component scissorCrossing_0;
	component doubleSwitch_0 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R5_command : in routeCommands := RELEASE;
			R6_command : in routeCommands := RELEASE;
			R69_command : in routeCommands := RELEASE;
			R70_command : in routeCommands := RELEASE;
			R77_command : in routeCommands := RELEASE;
			R78_command : in routeCommands := RELEASE;
			R79_command : in routeCommands := RELEASE;
			R80_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component doubleSwitch_0;
	component doubleSwitch_1 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			R36_command : in routeCommands := RELEASE;
			R37_command : in routeCommands := RELEASE;
			R65_command : in routeCommands := RELEASE;
			R66_command : in routeCommands := RELEASE;
			R82_command : in routeCommands := RELEASE;
			R83_command : in routeCommands := RELEASE;
			R89_command : in routeCommands := RELEASE;
			R90_command : in routeCommands := RELEASE;
			indication : in hex_char;
			command : out hex_char;
			correspondence : out hex_char
		);
	end component doubleSwitch_1;
	component railwaySignal_0 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R39_command : in routeCommands;
			--Ocupation level 0
			track_ne1 : in hex_char;
			correspondence_T01 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_0;
	component railwaySignal_1 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R1_command : in routeCommands;
			--Ocupation level 0
			track_ne1 : in hex_char;
			correspondence_T02 : out hex_char;
			correspondence_C78 : in hex_char;
			--Ocupation level 2
			track_ne9 : in hex_char;
			correspondence_J46 : in hex_char;
			s68W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_1;
	component railwaySignal_2 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R38_command : in routeCommands;
			R1_command : in routeCommands;
			--Ocupation level 0
			track_ne1 : in hex_char;
			correspondence_C78 : out hex_char;
			--Ocupation level 1
			track_ne9 : in hex_char;
			correspondence_J46 : in hex_char;
			s68W02_state : in hex_char;
			--Ocupation level 2
			track_ne95 : in hex_char;
			correspondence_L35 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_2;
	component railwaySignal_3 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R32_command : in routeCommands;
			--Ocupation level 0
			track_ne4 : in hex_char;
			correspondence_T03 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_3;
	component railwaySignal_4 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R10_command : in routeCommands;
			--Ocupation level 0
			track_ne4 : in hex_char;
			correspondence_L25 : out hex_char;
			--Ocupation level 1
			track_ne106 : in hex_char;
			correspondence_L42 : in hex_char;
			--Ocupation level 2
			track_ne99 : in hex_char;
			correspondence_P68 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_4;
	component railwaySignal_5 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R40_command : in routeCommands;
			--Ocupation level 0
			track_ne7 : in hex_char;
			correspondence_T05 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_5;
	component railwaySignal_6 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R2_command : in routeCommands;
			--Ocupation level 0
			track_ne7 : in hex_char;
			correspondence_T06 : out hex_char;
			correspondence_J43 : in hex_char;
			--Ocupation level 2
			track_ne9 : in hex_char;
			correspondence_J46 : in hex_char;
			s68W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_6;
	component railwaySignal_7 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R23_command : in routeCommands;
			R2_command : in routeCommands;
			--Ocupation level 0
			track_ne7 : in hex_char;
			correspondence_J43 : out hex_char;
			--Ocupation level 1
			track_ne9 : in hex_char;
			correspondence_J46 : in hex_char;
			s68W02_state : in hex_char;
			--Ocupation level 2
			track_ne95 : in hex_char;
			correspondence_L35 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_7;
	component railwaySignal_8 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R24_command : in routeCommands;
			R23_command : in routeCommands;
			R38_command : in routeCommands;
			--Ocupation level 0
			track_ne9 : in hex_char;
			correspondence_J46 : out hex_char;
			--Ocupation level 1
			track_ne95 : in hex_char;
			correspondence_L35 : in hex_char;
			correspondence_X50 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_8;
	component railwaySignal_9 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			R26_command : in routeCommands;
			--Ocupation level 0
			track_ne9 : in hex_char;
			correspondence_S80 : out hex_char;
			--Ocupation level 1
			track_ne1 : in hex_char;
			track_ne7 : in hex_char;
			correspondence_T01 : in hex_char;
			correspondence_T05 : in hex_char;
			s68W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_9;
	component railwaySignal_10 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R45_command : in routeCommands;
			--Ocupation level 0
			track_ne14 : in hex_char;
			correspondence_T07 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_10;
	component railwaySignal_11 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R3_command : in routeCommands;
			--Ocupation level 0
			track_ne14 : in hex_char;
			correspondence_T08 : out hex_char;
			--Ocupation level 1
			track_ne52 : in hex_char;
			correspondence_S146 : in hex_char;
			s69W04_state : in hex_char;
			--Ocupation level 2
			track_ne77 : in hex_char;
			correspondence_B145 : in hex_char;
			Sw03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_11;
	component railwaySignal_12 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R41_command : in routeCommands;
			R64_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne17 : in hex_char;
			correspondence_C82 : out hex_char;
			--Ocupation level 1
			track_ne59 : in hex_char;
			track_ne95 : in hex_char;
			correspondence_X51 : in hex_char;
			s69W03_state : in hex_char;
			--Ocupation level 2
			track_ne9 : in hex_char;
			correspondence_S80 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_12;
	component railwaySignal_13 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R63_command : in routeCommands;
			R43_command : in routeCommands;
			--Ocupation level 0
			track_ne17 : in hex_char;
			correspondence_C109 : out hex_char;
			--Ocupation level 1
			track_ne78 : in hex_char;
			correspondence_L33 : in hex_char;
			Sw06_state : in hex_char;
			--Ocupation level 2
			track_ne93 : in hex_char;
			correspondence_L34 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_13;
	component railwaySignal_14 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R27_command : in routeCommands;
			R47_command : in routeCommands;
			--Ocupation level 0
			track_ne23 : in hex_char;
			correspondence_P60 : out hex_char;
			--Ocupation level 1
			track_ne26 : in hex_char;
			correspondence_L27 : in hex_char;
			s70W02_state : in hex_char;
			--Ocupation level 2
			track_ne65 : in hex_char;
			correspondence_L30 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_14;
	component railwaySignal_15 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R46_command : in routeCommands;
			R50_command : in routeCommands;
			--Ocupation level 0
			track_ne23 : in hex_char;
			correspondence_B89 : out hex_char;
			--Ocupation level 1
			track_ne64 : in hex_char;
			track_ne103 : in hex_char;
			track_ne67 : in hex_char;
			correspondence_P64 : in hex_char;
			--Ocupation level 2
			track_ne70 : in hex_char;
			correspondence_L32 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_15;
	component railwaySignal_16 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R28_command : in routeCommands;
			R51_command : in routeCommands;
			--Ocupation level 0
			track_ne24 : in hex_char;
			correspondence_P63 : out hex_char;
			--Ocupation level 1
			track_ne64 : in hex_char;
			track_ne103 : in hex_char;
			track_ne67 : in hex_char;
			correspondence_P64 : in hex_char;
			--Ocupation level 2
			track_ne70 : in hex_char;
			correspondence_L32 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_16;
	component railwaySignal_17 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R49_command : in routeCommands;
			R48_command : in routeCommands;
			--Ocupation level 0
			track_ne24 : in hex_char;
			correspondence_B92 : out hex_char;
			--Ocupation level 1
			track_ne26 : in hex_char;
			correspondence_L27 : in hex_char;
			s70W02_state : in hex_char;
			--Ocupation level 2
			track_ne65 : in hex_char;
			correspondence_L30 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_17;
	component railwaySignal_18 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R11_command : in routeCommands;
			R27_command : in routeCommands;
			R49_command : in routeCommands;
			--Ocupation level 0
			track_ne26 : in hex_char;
			correspondence_L27 : out hex_char;
			--Ocupation level 1
			track_ne65 : in hex_char;
			correspondence_L30 : in hex_char;
			--Ocupation level 2
			track_ne102 : in hex_char;
			correspondence_C104 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_18;
	component railwaySignal_19 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R50_command : in routeCommands;
			R51_command : in routeCommands;
			R62_command : in routeCommands;
			--Ocupation level 0
			track_ne26 : in hex_char;
			correspondence_S93 : out hex_char;
			--Ocupation level 1
			track_ne23 : in hex_char;
			track_ne24 : in hex_char;
			correspondence_B89 : in hex_char;
			correspondence_P63 : in hex_char;
			s70W02_state : in hex_char;
			--Ocupation level 2
			track_ne67 : in hex_char;
			track_ne64 : in hex_char;
			track_ne103 : in hex_char;
			correspondence_P64 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_19;
	component railwaySignal_20 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R53_command : in routeCommands;
			R57_command : in routeCommands;
			--Ocupation level 0
			track_ne29 : in hex_char;
			correspondence_B96 : out hex_char;
			--Ocupation level 1
			track_ne30 : in hex_char;
			correspondence_S122 : in hex_char;
			Sw08_state : in hex_char;
			--Ocupation level 2
			track_ne87 : in hex_char;
			track_ne86 : in hex_char;
			track_ne91 : in hex_char;
			track_ne89 : in hex_char;
			track_ne90 : in hex_char;
			correspondence_T19 : in hex_char;
			correspondence_T15 : in hex_char;
			correspondence_T21 : in hex_char;
			Sw12_state : in hex_char;
			Sw11_state : in hex_char;
			Sw13_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_20;
	component railwaySignal_21 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R57_command : in routeCommands;
			R59_command : in routeCommands;
			--Ocupation level 0
			track_ne29 : in hex_char;
			correspondence_B101 : out hex_char;
			correspondence_B96 : in hex_char;
			--Ocupation level 2
			track_ne30 : in hex_char;
			correspondence_S122 : in hex_char;
			Sw08_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_21;
	component railwaySignal_22 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R54_command : in routeCommands;
			R55_command : in routeCommands;
			R7_command : in routeCommands;
			R8_command : in routeCommands;
			R73_command : in routeCommands;
			--Ocupation level 0
			track_ne30 : in hex_char;
			correspondence_S97 : out hex_char;
			--Ocupation level 1
			track_ne29 : in hex_char;
			track_ne110 : in hex_char;
			track_ne83 : in hex_char;
			correspondence_C138 : in hex_char;
			correspondence_C114 : in hex_char;
			Sw08_state : in hex_char;
			Sw09_state : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			track_ne101 : in hex_char;
			track_ne44 : in hex_char;
			track_ne32 : in hex_char;
			correspondence_S105 : in hex_char;
			correspondence_C100 : in hex_char;
			Sw41_state : in hex_char;
			Sw04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_22;
	component railwaySignal_23 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			R52_command : in routeCommands;
			R53_command : in routeCommands;
			--Ocupation level 0
			track_ne30 : in hex_char;
			correspondence_S122 : out hex_char;
			--Ocupation level 1
			track_ne89 : in hex_char;
			track_ne91 : in hex_char;
			track_ne87 : in hex_char;
			track_ne86 : in hex_char;
			track_ne90 : in hex_char;
			correspondence_T19 : in hex_char;
			correspondence_T15 : in hex_char;
			correspondence_T21 : in hex_char;
			Sw12_state : in hex_char;
			Sw11_state : in hex_char;
			Sw13_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_23;
	component railwaySignal_24 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R56_command : in routeCommands;
			R5_command : in routeCommands;
			R67_command : in routeCommands;
			R77_command : in routeCommands;
			--Ocupation level 0
			track_ne32 : in hex_char;
			correspondence_C100 : out hex_char;
			--Ocupation level 1
			track_ne110 : in hex_char;
			correspondence_C138 : in hex_char;
			Sw09_state : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			track_ne101 : in hex_char;
			track_ne44 : in hex_char;
			correspondence_S105 : in hex_char;
			Sw41_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_24;
	component railwaySignal_25 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R58_command : in routeCommands;
			--Ocupation level 0
			track_ne32 : in hex_char;
			correspondence_S115 : out hex_char;
			--Ocupation level 1
			track_ne83 : in hex_char;
			track_ne82 : in hex_char;
			track_ne41 : in hex_char;
			track_ne84 : in hex_char;
			correspondence_C95 : in hex_char;
			correspondence_P58 : in hex_char;
			correspondence_T13 : in hex_char;
			Sw04_state : in hex_char;
			Sw05_state : in hex_char;
			--Ocupation level 2
			track_ne30 : in hex_char;
			correspondence_S122 : in hex_char;
			Sw08_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_25;
	component railwaySignal_26 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R69_command : in routeCommands;
			R79_command : in routeCommands;
			--Ocupation level 0
			track_ne41 : in hex_char;
			correspondence_P58 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_26;
	component railwaySignal_27 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			--Ocupation level 0
			track_ne41 : in hex_char;
			correspondence_B130 : out hex_char;
			--Ocupation level 1
			track_ne82 : in hex_char;
			track_ne32 : in hex_char;
			track_ne85 : in hex_char;
			track_ne100 : in hex_char;
			track_ne101 : in hex_char;
			track_ne44 : in hex_char;
			correspondence_C100 : in hex_char;
			correspondence_S105 : in hex_char;
			Sw04_state : in hex_char;
			Sw05_state : in hex_char;
			Sw41_state : in hex_char;
			--Ocupation level 2
			track_ne110 : in hex_char;
			track_ne26 : in hex_char;
			track_ne43 : in hex_char;
			track_ne102 : in hex_char;
			track_ne48 : in hex_char;
			track_ne65 : in hex_char;
			correspondence_C138 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_S93 : in hex_char;
			Sw09_state : in hex_char;
			s71W01_state : in hex_char;
			s71W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_27;
	component railwaySignal_28 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R12_command : in routeCommands;
			R60_command : in routeCommands;
			--Ocupation level 0
			track_ne44 : in hex_char;
			correspondence_L28 : out hex_char;
			--Ocupation level 1
			track_ne101 : in hex_char;
			correspondence_L40 : in hex_char;
			--Ocupation level 2
			track_ne100 : in hex_char;
			correspondence_S139 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_28;
	component railwaySignal_29 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			R6_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			--Ocupation level 0
			track_ne44 : in hex_char;
			correspondence_S105 : out hex_char;
			--Ocupation level 1
			track_ne43 : in hex_char;
			track_ne48 : in hex_char;
			track_ne102 : in hex_char;
			track_ne65 : in hex_char;
			track_ne26 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_S93 : in hex_char;
			s71W01_state : in hex_char;
			s71W02_state : in hex_char;
			--Ocupation level 2
			track_ne23 : in hex_char;
			track_ne24 : in hex_char;
			correspondence_B89 : in hex_char;
			correspondence_P63 : in hex_char;
			s70W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_29;
	component railwaySignal_30 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			--Ocupation level 0
			track_ne47 : in hex_char;
			correspondence_T11 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_30;
	component railwaySignal_31 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			--Ocupation level 0
			track_ne47 : in hex_char;
			correspondence_T12 : out hex_char;
			--Ocupation level 1
			track_ne48 : in hex_char;
			correspondence_L29 : in hex_char;
			s71W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_31;
	component railwaySignal_32 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R4_command : in routeCommands;
			R61_command : in routeCommands;
			--Ocupation level 0
			track_ne48 : in hex_char;
			correspondence_L29 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_32;
	component railwaySignal_33 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R42_command : in routeCommands;
			R43_command : in routeCommands;
			R25_command : in routeCommands;
			--Ocupation level 0
			track_ne59 : in hex_char;
			correspondence_S83 : out hex_char;
			--Ocupation level 1
			track_ne11 : in hex_char;
			track_ne52 : in hex_char;
			track_ne17 : in hex_char;
			correspondence_S146 : in hex_char;
			correspondence_C109 : in hex_char;
			s69W03_state : in hex_char;
			s69W04_state : in hex_char;
			--Ocupation level 2
			track_ne77 : in hex_char;
			track_ne78 : in hex_char;
			correspondence_B145 : in hex_char;
			correspondence_L33 : in hex_char;
			Sw03_state : in hex_char;
			Sw06_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_33;
	component railwaySignal_34 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R47_command : in routeCommands;
			R48_command : in routeCommands;
			R21_command : in routeCommands;
			--Ocupation level 0
			track_ne64 : in hex_char;
			correspondence_S90 : out hex_char;
			--Ocupation level 1
			track_ne23 : in hex_char;
			track_ne24 : in hex_char;
			correspondence_P60 : in hex_char;
			correspondence_B92 : in hex_char;
			s70W01_state : in hex_char;
			--Ocupation level 2
			track_ne26 : in hex_char;
			correspondence_L27 : in hex_char;
			s70W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_34;
	component railwaySignal_35 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R13_command : in routeCommands;
			R11_command : in routeCommands;
			--Ocupation level 0
			track_ne65 : in hex_char;
			correspondence_L30 : out hex_char;
			--Ocupation level 1
			track_ne102 : in hex_char;
			correspondence_C104 : in hex_char;
			--Ocupation level 2
			track_ne44 : in hex_char;
			correspondence_L28 : in hex_char;
			s71W01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_35;
	component railwaySignal_36 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R29_command : in routeCommands;
			R28_command : in routeCommands;
			R46_command : in routeCommands;
			--Ocupation level 0
			track_ne67 : in hex_char;
			correspondence_P64 : out hex_char;
			--Ocupation level 1
			track_ne70 : in hex_char;
			correspondence_L32 : in hex_char;
			--Ocupation level 2
			track_ne104 : in hex_char;
			track_ne21 : in hex_char;
			correspondence_P73 : in hex_char;
			Sw03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_36;
	component railwaySignal_37 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R30_command : in routeCommands;
			--Ocupation level 0
			track_ne67 : in hex_char;
			correspondence_P65 : out hex_char;
			--Ocupation level 1
			track_ne103 : in hex_char;
			correspondence_L41 : in hex_char;
			--Ocupation level 2
			track_ne64 : in hex_char;
			correspondence_S90 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_37;
	component railwaySignal_38 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R14_command : in routeCommands;
			R29_command : in routeCommands;
			R87_command : in routeCommands;
			--Ocupation level 0
			track_ne70 : in hex_char;
			correspondence_L32 : out hex_char;
			--Ocupation level 1
			track_ne104 : in hex_char;
			track_ne21 : in hex_char;
			correspondence_P73 : in hex_char;
			Sw03_state : in hex_char;
			--Ocupation level 2
			track_ne97 : in hex_char;
			track_ne94 : in hex_char;
			track_ne79 : in hex_char;
			track_ne78 : in hex_char;
			track_ne99 : in hex_char;
			correspondence_L33 : in hex_char;
			correspondence_P69 : in hex_char;
			Sw06_state : in hex_char;
			Sw07_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_38;
	component railwaySignal_39 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R15_command : in routeCommands;
			R36_command : in routeCommands;
			R63_command : in routeCommands;
			R89_command : in routeCommands;
			--Ocupation level 0
			track_ne78 : in hex_char;
			correspondence_L33 : out hex_char;
			--Ocupation level 1
			track_ne93 : in hex_char;
			correspondence_L34 : in hex_char;
			--Ocupation level 2
			track_ne96 : in hex_char;
			correspondence_P71 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_39;
	component railwaySignal_40 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R64_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R33_command : in routeCommands;
			--Ocupation level 0
			track_ne78 : in hex_char;
			correspondence_S110 : out hex_char;
			--Ocupation level 1
			track_ne17 : in hex_char;
			track_ne79 : in hex_char;
			track_ne77 : in hex_char;
			track_ne21 : in hex_char;
			correspondence_C82 : in hex_char;
			correspondence_B133 : in hex_char;
			correspondence_P72 : in hex_char;
			Sw06_state : in hex_char;
			Sw07_state : in hex_char;
			--Ocupation level 2
			track_ne59 : in hex_char;
			track_ne95 : in hex_char;
			track_ne52 : in hex_char;
			correspondence_X51 : in hex_char;
			correspondence_S86 : in hex_char;
			correspondence_S144 : in hex_char;
			s69W03_state : in hex_char;
			Sw03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_40;
	component railwaySignal_41 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R52_command : in routeCommands;
			R68_command : in routeCommands;
			--Ocupation level 0
			track_ne83 : in hex_char;
			correspondence_C95 : out hex_char;
			--Ocupation level 1
			track_ne30 : in hex_char;
			correspondence_S122 : in hex_char;
			Sw08_state : in hex_char;
			--Ocupation level 2
			track_ne87 : in hex_char;
			track_ne86 : in hex_char;
			track_ne91 : in hex_char;
			track_ne89 : in hex_char;
			track_ne90 : in hex_char;
			correspondence_T19 : in hex_char;
			correspondence_T15 : in hex_char;
			correspondence_T21 : in hex_char;
			Sw12_state : in hex_char;
			Sw11_state : in hex_char;
			Sw13_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_41;
	component railwaySignal_42 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R67_command : in routeCommands;
			R55_command : in routeCommands;
			--Ocupation level 0
			track_ne83 : in hex_char;
			correspondence_C114 : out hex_char;
			--Ocupation level 1
			track_ne32 : in hex_char;
			correspondence_C100 : in hex_char;
			Sw04_state : in hex_char;
			--Ocupation level 2
			track_ne110 : in hex_char;
			correspondence_C138 : in hex_char;
			Sw09_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_42;
	component railwaySignal_43 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R70_command : in routeCommands;
			R80_command : in routeCommands;
			--Ocupation level 0
			track_ne84 : in hex_char;
			correspondence_T13 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_43;
	component railwaySignal_44 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R5_command : in routeCommands;
			R6_command : in routeCommands;
			--Ocupation level 0
			track_ne84 : in hex_char;
			correspondence_T14 : out hex_char;
			--Ocupation level 1
			track_ne82 : in hex_char;
			track_ne32 : in hex_char;
			track_ne85 : in hex_char;
			track_ne100 : in hex_char;
			track_ne101 : in hex_char;
			track_ne44 : in hex_char;
			correspondence_C100 : in hex_char;
			correspondence_S105 : in hex_char;
			Sw04_state : in hex_char;
			Sw05_state : in hex_char;
			Sw41_state : in hex_char;
			--Ocupation level 2
			track_ne110 : in hex_char;
			track_ne26 : in hex_char;
			track_ne43 : in hex_char;
			track_ne102 : in hex_char;
			track_ne48 : in hex_char;
			track_ne65 : in hex_char;
			correspondence_C138 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_S93 : in hex_char;
			Sw09_state : in hex_char;
			s71W01_state : in hex_char;
			s71W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_44;
	component railwaySignal_45 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R71_command : in routeCommands;
			R75_command : in routeCommands;
			--Ocupation level 0
			track_ne86 : in hex_char;
			correspondence_T15 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_45;
	component railwaySignal_46 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R72_command : in routeCommands;
			R73_command : in routeCommands;
			--Ocupation level 0
			track_ne86 : in hex_char;
			correspondence_S119 : out hex_char;
			--Ocupation level 1
			track_ne88 : in hex_char;
			track_ne87 : in hex_char;
			track_ne91 : in hex_char;
			track_ne30 : in hex_char;
			correspondence_T17 : in hex_char;
			correspondence_S97 : in hex_char;
			Sw11_state : in hex_char;
			Sw12_state : in hex_char;
			Sw13_state : in hex_char;
			--Ocupation level 2
			track_ne83 : in hex_char;
			track_ne29 : in hex_char;
			track_ne110 : in hex_char;
			correspondence_C138 : in hex_char;
			correspondence_C114 : in hex_char;
			Sw08_state : in hex_char;
			Sw09_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_46;
	component railwaySignal_47 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R72_command : in routeCommands;
			--Ocupation level 0
			track_ne88 : in hex_char;
			correspondence_T17 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_47;
	component railwaySignal_48 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R71_command : in routeCommands;
			--Ocupation level 0
			track_ne88 : in hex_char;
			correspondence_C118 : out hex_char;
			--Ocupation level 1
			track_ne86 : in hex_char;
			correspondence_T15 : in hex_char;
			Sw11_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_48;
	component railwaySignal_49 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R74_command : in routeCommands;
			--Ocupation level 0
			track_ne89 : in hex_char;
			correspondence_T19 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_49;
	component railwaySignal_50 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R7_command : in routeCommands;
			--Ocupation level 0
			track_ne89 : in hex_char;
			correspondence_T20 : out hex_char;
			--Ocupation level 1
			track_ne30 : in hex_char;
			correspondence_S97 : in hex_char;
			Sw12_state : in hex_char;
			--Ocupation level 2
			track_ne83 : in hex_char;
			track_ne29 : in hex_char;
			track_ne110 : in hex_char;
			correspondence_C138 : in hex_char;
			correspondence_C114 : in hex_char;
			Sw08_state : in hex_char;
			Sw09_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_50;
	component railwaySignal_51 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R76_command : in routeCommands;
			--Ocupation level 0
			track_ne90 : in hex_char;
			correspondence_T21 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_51;
	component railwaySignal_52 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R8_command : in routeCommands;
			--Ocupation level 0
			track_ne90 : in hex_char;
			correspondence_T22 : out hex_char;
			--Ocupation level 1
			track_ne91 : in hex_char;
			track_ne30 : in hex_char;
			correspondence_S97 : in hex_char;
			Sw12_state : in hex_char;
			Sw13_state : in hex_char;
			--Ocupation level 2
			track_ne83 : in hex_char;
			track_ne29 : in hex_char;
			track_ne110 : in hex_char;
			correspondence_C138 : in hex_char;
			correspondence_C114 : in hex_char;
			Sw08_state : in hex_char;
			Sw09_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_52;
	component railwaySignal_53 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R16_command : in routeCommands;
			R15_command : in routeCommands;
			--Ocupation level 0
			track_ne93 : in hex_char;
			correspondence_L34 : out hex_char;
			--Ocupation level 1
			track_ne96 : in hex_char;
			correspondence_P71 : in hex_char;
			--Ocupation level 2
			track_ne98 : in hex_char;
			correspondence_L38 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_53;
	component railwaySignal_54 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			R18_command : in routeCommands;
			--Ocupation level 0
			track_ne94 : in hex_char;
			correspondence_S135 : out hex_char;
			--Ocupation level 1
			track_ne77 : in hex_char;
			track_ne21 : in hex_char;
			correspondence_B133 : in hex_char;
			correspondence_P72 : in hex_char;
			Sw07_state : in hex_char;
			--Ocupation level 2
			track_ne52 : in hex_char;
			correspondence_S86 : in hex_char;
			correspondence_S144 : in hex_char;
			Sw03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_54;
	component railwaySignal_55 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R17_command : in routeCommands;
			R24_command : in routeCommands;
			--Ocupation level 0
			track_ne95 : in hex_char;
			correspondence_L35 : out hex_char;
			correspondence_X50 : in hex_char;
			--Ocupation level 2
			track_ne59 : in hex_char;
			correspondence_S83 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_55;
	component railwaySignal_56 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R25_command : in routeCommands;
			R17_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne95 : in hex_char;
			correspondence_X50 : out hex_char;
			--Ocupation level 1
			track_ne59 : in hex_char;
			correspondence_S83 : in hex_char;
			--Ocupation level 2
			track_ne17 : in hex_char;
			track_ne11 : in hex_char;
			track_ne52 : in hex_char;
			correspondence_S146 : in hex_char;
			correspondence_C109 : in hex_char;
			s69W03_state : in hex_char;
			s69W04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_56;
	component railwaySignal_57 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R26_command : in routeCommands;
			R41_command : in routeCommands;
			R44_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne95 : in hex_char;
			correspondence_X51 : out hex_char;
			--Ocupation level 1
			track_ne9 : in hex_char;
			correspondence_S80 : in hex_char;
			--Ocupation level 2
			track_ne7 : in hex_char;
			track_ne1 : in hex_char;
			correspondence_T01 : in hex_char;
			correspondence_T05 : in hex_char;
			s68W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_57;
	component railwaySignal_58 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R33_command : in routeCommands;
			R9_command : in routeCommands;
			--Ocupation level 0
			track_ne96 : in hex_char;
			correspondence_P70 : out hex_char;
			--Ocupation level 1
			track_ne93 : in hex_char;
			track_ne78 : in hex_char;
			correspondence_S110 : in hex_char;
			--Ocupation level 2
			track_ne17 : in hex_char;
			track_ne79 : in hex_char;
			track_ne21 : in hex_char;
			track_ne77 : in hex_char;
			correspondence_C82 : in hex_char;
			correspondence_B133 : in hex_char;
			correspondence_P72 : in hex_char;
			Sw06_state : in hex_char;
			Sw07_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_58;
	component railwaySignal_59 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R34_command : in routeCommands;
			R16_command : in routeCommands;
			--Ocupation level 0
			track_ne96 : in hex_char;
			correspondence_P71 : out hex_char;
			--Ocupation level 1
			track_ne98 : in hex_char;
			correspondence_L38 : in hex_char;
			--Ocupation level 2
			track_ne105 : in hex_char;
			correspondence_T23 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_59;
	component railwaySignal_60 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R18_command : in routeCommands;
			R31_command : in routeCommands;
			--Ocupation level 0
			track_ne97 : in hex_char;
			correspondence_L37 : out hex_char;
			--Ocupation level 1
			track_ne94 : in hex_char;
			correspondence_S135 : in hex_char;
			--Ocupation level 2
			track_ne21 : in hex_char;
			track_ne77 : in hex_char;
			correspondence_B133 : in hex_char;
			correspondence_P72 : in hex_char;
			Sw07_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_60;
	component railwaySignal_61 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R19_command : in routeCommands;
			R34_command : in routeCommands;
			--Ocupation level 0
			track_ne98 : in hex_char;
			correspondence_L38 : out hex_char;
			--Ocupation level 1
			track_ne105 : in hex_char;
			correspondence_T23 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_61;
	component railwaySignal_62 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R31_command : in routeCommands;
			R22_command : in routeCommands;
			--Ocupation level 0
			track_ne99 : in hex_char;
			correspondence_P68 : out hex_char;
			--Ocupation level 1
			track_ne97 : in hex_char;
			correspondence_L37 : in hex_char;
			--Ocupation level 2
			track_ne94 : in hex_char;
			correspondence_S135 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_62;
	component railwaySignal_63 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R32_command : in routeCommands;
			R37_command : in routeCommands;
			R90_command : in routeCommands;
			--Ocupation level 0
			track_ne99 : in hex_char;
			correspondence_P69 : out hex_char;
			--Ocupation level 1
			track_ne106 : in hex_char;
			track_ne4 : in hex_char;
			correspondence_T03 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_63;
	component railwaySignal_64 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			R20_command : in routeCommands;
			--Ocupation level 0
			track_ne100 : in hex_char;
			correspondence_S139 : out hex_char;
			--Ocupation level 1
			track_ne110 : in hex_char;
			track_ne85 : in hex_char;
			correspondence_S102 : in hex_char;
			correspondence_S131 : in hex_char;
			Sw41_state : in hex_char;
			--Ocupation level 2
			track_ne32 : in hex_char;
			track_ne29 : in hex_char;
			track_ne84 : in hex_char;
			track_ne41 : in hex_char;
			correspondence_S115 : in hex_char;
			correspondence_B101 : in hex_char;
			correspondence_P58 : in hex_char;
			correspondence_T13 : in hex_char;
			Sw09_state : in hex_char;
			Sw05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_64;
	component railwaySignal_65 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R20_command : in routeCommands;
			R12_command : in routeCommands;
			--Ocupation level 0
			track_ne101 : in hex_char;
			correspondence_L40 : out hex_char;
			--Ocupation level 1
			track_ne100 : in hex_char;
			correspondence_S139 : in hex_char;
			--Ocupation level 2
			track_ne85 : in hex_char;
			track_ne110 : in hex_char;
			correspondence_S102 : in hex_char;
			correspondence_S131 : in hex_char;
			Sw41_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_65;
	component railwaySignal_66 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R60_command : in routeCommands;
			R13_command : in routeCommands;
			--Ocupation level 0
			track_ne102 : in hex_char;
			correspondence_C104 : out hex_char;
			--Ocupation level 1
			track_ne44 : in hex_char;
			correspondence_L28 : in hex_char;
			s71W01_state : in hex_char;
			--Ocupation level 2
			track_ne101 : in hex_char;
			correspondence_L40 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_66;
	component railwaySignal_67 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R21_command : in routeCommands;
			R30_command : in routeCommands;
			--Ocupation level 0
			track_ne103 : in hex_char;
			correspondence_L41 : out hex_char;
			--Ocupation level 1
			track_ne64 : in hex_char;
			correspondence_S90 : in hex_char;
			--Ocupation level 2
			track_ne23 : in hex_char;
			track_ne24 : in hex_char;
			correspondence_P60 : in hex_char;
			correspondence_B92 : in hex_char;
			s70W01_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_67;
	component railwaySignal_68 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R19_command : in routeCommands;
			--Ocupation level 0
			track_ne105 : in hex_char;
			correspondence_T23 : out hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_68;
	component railwaySignal_69 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R9_command : in routeCommands;
			--Ocupation level 0
			track_ne105 : in hex_char;
			correspondence_T24 : out hex_char;
			--Ocupation level 1
			track_ne98 : in hex_char;
			track_ne96 : in hex_char;
			correspondence_P70 : in hex_char;
			--Ocupation level 2
			track_ne93 : in hex_char;
			track_ne78 : in hex_char;
			correspondence_S110 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_69;
	component railwaySignal_70 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R22_command : in routeCommands;
			R10_command : in routeCommands;
			--Ocupation level 0
			track_ne106 : in hex_char;
			correspondence_L42 : out hex_char;
			--Ocupation level 1
			track_ne99 : in hex_char;
			correspondence_P68 : in hex_char;
			--Ocupation level 2
			track_ne97 : in hex_char;
			correspondence_L37 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_70;
	component railwaySignal_71 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			R86_command : in routeCommands;
			--Ocupation level 0
			track_ne85 : in hex_char;
			correspondence_S131 : out hex_char;
			--Ocupation level 1
			track_ne41 : in hex_char;
			track_ne84 : in hex_char;
			correspondence_P58 : in hex_char;
			correspondence_T13 : in hex_char;
			Sw05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_71;
	component railwaySignal_72 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R81_command : in routeCommands;
			R65_command : in routeCommands;
			R82_command : in routeCommands;
			--Ocupation level 0
			track_ne77 : in hex_char;
			correspondence_B133 : out hex_char;
			--Ocupation level 1
			track_ne52 : in hex_char;
			correspondence_S86 : in hex_char;
			Sw03_state : in hex_char;
			--Ocupation level 2
			track_ne59 : in hex_char;
			track_ne11 : in hex_char;
			track_ne14 : in hex_char;
			track_ne95 : in hex_char;
			correspondence_X51 : in hex_char;
			correspondence_T07 : in hex_char;
			s69W03_state : in hex_char;
			s69W04_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_72;
	component railwaySignal_73 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R89_command : in routeCommands;
			R90_command : in routeCommands;
			R91_command : in routeCommands;
			--Ocupation level 0
			track_ne77 : in hex_char;
			correspondence_B145 : out hex_char;
			--Ocupation level 1
			track_ne79 : in hex_char;
			track_ne78 : in hex_char;
			track_ne94 : in hex_char;
			track_ne97 : in hex_char;
			track_ne99 : in hex_char;
			correspondence_L33 : in hex_char;
			correspondence_P69 : in hex_char;
			Sw06_state : in hex_char;
			Sw07_state : in hex_char;
			--Ocupation level 2
			track_ne93 : in hex_char;
			track_ne4 : in hex_char;
			track_ne106 : in hex_char;
			correspondence_L34 : in hex_char;
			correspondence_T03 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_73;
	component railwaySignal_74 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			--Ocupation level 0
			track_ne104 : in hex_char;
			correspondence_B143 : out hex_char;
			--Ocupation level 1
			track_ne70 : in hex_char;
			correspondence_L32 : in hex_char;
			--Ocupation level 2
			track_ne21 : in hex_char;
			correspondence_P73 : in hex_char;
			Sw03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_74;
	component railwaySignal_75 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R44_command : in routeCommands;
			R45_command : in routeCommands;
			R81_command : in routeCommands;
			Lc01_state : in hex_char;
			--Ocupation level 0
			track_ne52 : in hex_char;
			correspondence_S86 : out hex_char;
			--Ocupation level 1
			track_ne11 : in hex_char;
			track_ne59 : in hex_char;
			track_ne95 : in hex_char;
			track_ne14 : in hex_char;
			correspondence_X51 : in hex_char;
			correspondence_T07 : in hex_char;
			s69W03_state : in hex_char;
			s69W04_state : in hex_char;
			--Ocupation level 2
			track_ne9 : in hex_char;
			correspondence_S80 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_75;
	component railwaySignal_76 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R91_command : in routeCommands;
			R3_command : in routeCommands;
			R42_command : in routeCommands;
			--Ocupation level 0
			track_ne52 : in hex_char;
			correspondence_S146 : out hex_char;
			--Ocupation level 1
			track_ne77 : in hex_char;
			correspondence_B145 : in hex_char;
			Sw03_state : in hex_char;
			--Ocupation level 2
			track_ne97 : in hex_char;
			track_ne94 : in hex_char;
			track_ne79 : in hex_char;
			track_ne78 : in hex_char;
			track_ne99 : in hex_char;
			correspondence_L33 : in hex_char;
			correspondence_P69 : in hex_char;
			Sw06_state : in hex_char;
			Sw07_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_76;
	component railwaySignal_77 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R35_command : in routeCommands;
			R66_command : in routeCommands;
			R83_command : in routeCommands;
			--Ocupation level 0
			track_ne21 : in hex_char;
			correspondence_P72 : out hex_char;
			correspondence_S144 : in hex_char;
			--Ocupation level 2
			track_ne104 : in hex_char;
			correspondence_B143 : in hex_char;
			Sw03_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_77;
	component railwaySignal_78 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R36_command : in routeCommands;
			R37_command : in routeCommands;
			R14_command : in routeCommands;
			--Ocupation level 0
			track_ne21 : in hex_char;
			correspondence_P73 : out hex_char;
			--Ocupation level 1
			track_ne79 : in hex_char;
			track_ne78 : in hex_char;
			track_ne94 : in hex_char;
			track_ne97 : in hex_char;
			track_ne99 : in hex_char;
			correspondence_L33 : in hex_char;
			correspondence_P69 : in hex_char;
			Sw06_state : in hex_char;
			Sw07_state : in hex_char;
			--Ocupation level 2
			track_ne93 : in hex_char;
			track_ne4 : in hex_char;
			track_ne106 : in hex_char;
			correspondence_L34 : in hex_char;
			correspondence_T03 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_78;
	component railwaySignal_79 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R88_command : in routeCommands;
			R35_command : in routeCommands;
			--Ocupation level 0
			track_ne21 : in hex_char;
			correspondence_S144 : out hex_char;
			--Ocupation level 1
			track_ne104 : in hex_char;
			correspondence_B143 : in hex_char;
			Sw03_state : in hex_char;
			--Ocupation level 2
			track_ne70 : in hex_char;
			correspondence_L32 : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_79;
	component railwaySignal_80 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R58_command : in routeCommands;
			R59_command : in routeCommands;
			R85_command : in routeCommands;
			--Ocupation level 0
			track_ne110 : in hex_char;
			correspondence_S102 : out hex_char;
			--Ocupation level 1
			track_ne32 : in hex_char;
			track_ne29 : in hex_char;
			correspondence_S115 : in hex_char;
			correspondence_B101 : in hex_char;
			Sw09_state : in hex_char;
			--Ocupation level 2
			track_ne84 : in hex_char;
			track_ne83 : in hex_char;
			track_ne41 : in hex_char;
			track_ne82 : in hex_char;
			correspondence_C95 : in hex_char;
			correspondence_P58 : in hex_char;
			correspondence_T13 : in hex_char;
			correspondence_B96 : in hex_char;
			Sw04_state : in hex_char;
			Sw05_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_80;
	component railwaySignal_81 is
		port(
			clock : in std_logic;
			reset : in std_logic;
			R84_command : in routeCommands;
			R54_command : in routeCommands;
			R56_command : in routeCommands;
			--Ocupation level 0
			track_ne110 : in hex_char;
			correspondence_C138 : out hex_char;
			--Ocupation level 1
			track_ne100 : in hex_char;
			track_ne101 : in hex_char;
			track_ne44 : in hex_char;
			correspondence_S105 : in hex_char;
			Sw41_state : in hex_char;
			--Ocupation level 2
			track_ne26 : in hex_char;
			track_ne43 : in hex_char;
			track_ne102 : in hex_char;
			track_ne48 : in hex_char;
			track_ne65 : in hex_char;
			correspondence_L29 : in hex_char;
			correspondence_S93 : in hex_char;
			s71W01_state : in hex_char;
			s71W02_state : in hex_char;
			indication : in hex_char;
			command : out hex_char
		);
	end component railwaySignal_81;
	component node_0 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R1_command : in routeCommands;
			R38_command : in routeCommands;
			R39_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_0;
	component node_1 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R10_command : in routeCommands;
			R32_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_1;
	component node_2 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R2_command : in routeCommands;
			R23_command : in routeCommands;
			R40_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_2;
	component node_3 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R23_command : in routeCommands;
			R24_command : in routeCommands;
			R26_command : in routeCommands;
			R38_command : in routeCommands;
			R39_command : in routeCommands;
			R40_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_3;
	component node_4 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_4;
	component node_5 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R3_command : in routeCommands;
			R45_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_5;
	component node_6 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R41_command : in routeCommands;
			R43_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_6;
	component node_7 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R27_command : in routeCommands;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			R50_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_7;
	component node_8 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R28_command : in routeCommands;
			R48_command : in routeCommands;
			R49_command : in routeCommands;
			R51_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_8;
	component node_9 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R11_command : in routeCommands;
			R27_command : in routeCommands;
			R49_command : in routeCommands;
			R50_command : in routeCommands;
			R51_command : in routeCommands;
			R62_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_9;
	component node_10 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R57_command : in routeCommands;
			R59_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_10;
	component node_11 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R7_command : in routeCommands;
			R8_command : in routeCommands;
			R52_command : in routeCommands;
			R53_command : in routeCommands;
			R54_command : in routeCommands;
			R55_command : in routeCommands;
			R73_command : in routeCommands;
			R74_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_11;
	component node_12 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R5_command : in routeCommands;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R67_command : in routeCommands;
			R68_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R77_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_12;
	component node_13 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R69_command : in routeCommands;
			R77_command : in routeCommands;
			R78_command : in routeCommands;
			R79_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_13;
	component node_14 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R61_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_14;
	component node_15 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R6_command : in routeCommands;
			R12_command : in routeCommands;
			R60_command : in routeCommands;
			R61_command : in routeCommands;
			R62_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_15;
	component node_16 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R4_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_16;
	component node_17 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R4_command : in routeCommands;
			R61_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_17;
	component node_18 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R25_command : in routeCommands;
			R41_command : in routeCommands;
			R42_command : in routeCommands;
			R43_command : in routeCommands;
			R44_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_18;
	component node_19 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R21_command : in routeCommands;
			R28_command : in routeCommands;
			R46_command : in routeCommands;
			R47_command : in routeCommands;
			R48_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_19;
	component node_20 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R11_command : in routeCommands;
			R13_command : in routeCommands;
			R62_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_20;
	component node_21 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R28_command : in routeCommands;
			R29_command : in routeCommands;
			R30_command : in routeCommands;
			R46_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_21;
	component node_22 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R14_command : in routeCommands;
			R29_command : in routeCommands;
			R87_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_22;
	component node_23 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R15_command : in routeCommands;
			R33_command : in routeCommands;
			R36_command : in routeCommands;
			R63_command : in routeCommands;
			R64_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R89_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_23;
	component node_24 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R36_command : in routeCommands;
			R65_command : in routeCommands;
			R66_command : in routeCommands;
			R89_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_24;
	component node_25 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R5_command : in routeCommands;
			R69_command : in routeCommands;
			R70_command : in routeCommands;
			R77_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_25;
	component node_26 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R52_command : in routeCommands;
			R55_command : in routeCommands;
			R67_command : in routeCommands;
			R68_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_26;
	component node_27 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R5_command : in routeCommands;
			R6_command : in routeCommands;
			R70_command : in routeCommands;
			R80_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_27;
	component node_28 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_28;
	component node_29 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_29;
	component node_30 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R71_command : in routeCommands;
			R72_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_30;
	component node_31 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R7_command : in routeCommands;
			R74_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_31;
	component node_32 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R8_command : in routeCommands;
			R76_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_32;
	component node_33 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R8_command : in routeCommands;
			R73_command : in routeCommands;
			R75_command : in routeCommands;
			R76_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_33;
	component node_34 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R15_command : in routeCommands;
			R16_command : in routeCommands;
			R33_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_34;
	component node_35 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R18_command : in routeCommands;
			R37_command : in routeCommands;
			R82_command : in routeCommands;
			R83_command : in routeCommands;
			R90_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_35;
	component node_36 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R17_command : in routeCommands;
			R24_command : in routeCommands;
			R25_command : in routeCommands;
			R26_command : in routeCommands;
			R41_command : in routeCommands;
			R44_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_36;
	component node_37 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R9_command : in routeCommands;
			R16_command : in routeCommands;
			R33_command : in routeCommands;
			R34_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_37;
	component node_38 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R18_command : in routeCommands;
			R31_command : in routeCommands;
			R37_command : in routeCommands;
			R90_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_38;
	component node_39 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R9_command : in routeCommands;
			R19_command : in routeCommands;
			R34_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_39;
	component node_40 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R22_command : in routeCommands;
			R31_command : in routeCommands;
			R32_command : in routeCommands;
			R37_command : in routeCommands;
			R90_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_40;
	component node_41 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R6_command : in routeCommands;
			R20_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			R86_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_41;
	component node_42 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R6_command : in routeCommands;
			R12_command : in routeCommands;
			R20_command : in routeCommands;
			R78_command : in routeCommands;
			R84_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_42;
	component node_43 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R13_command : in routeCommands;
			R60_command : in routeCommands;
			R62_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_43;
	component node_44 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R21_command : in routeCommands;
			R28_command : in routeCommands;
			R30_command : in routeCommands;
			R46_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_44;
	component node_45 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R9_command : in routeCommands;
			R19_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_45;
	component node_46 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R10_command : in routeCommands;
			R22_command : in routeCommands;
			R32_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_46;
	component node_47 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R6_command : in routeCommands;
			R78_command : in routeCommands;
			R79_command : in routeCommands;
			R80_command : in routeCommands;
			R86_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_47;
	component node_48 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R65_command : in routeCommands;
			R81_command : in routeCommands;
			R82_command : in routeCommands;
			R89_command : in routeCommands;
			R90_command : in routeCommands;
			R91_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_48;
	component node_49 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R14_command : in routeCommands;
			R87_command : in routeCommands;
			R88_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_49;
	component node_50 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R3_command : in routeCommands;
			R42_command : in routeCommands;
			R44_command : in routeCommands;
			R45_command : in routeCommands;
			R81_command : in routeCommands;
			R91_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_50;
	component node_51 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R14_command : in routeCommands;
			R35_command : in routeCommands;
			R36_command : in routeCommands;
			R37_command : in routeCommands;
			R66_command : in routeCommands;
			R83_command : in routeCommands;
			R88_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_51;
	component node_52 is
		port(
			reset : in std_logic;
			track_i : in hex_char;
			R54_command : in routeCommands;
			R56_command : in routeCommands;
			R58_command : in routeCommands;
			R59_command : in routeCommands;
			R84_command : in routeCommands;
			R85_command : in routeCommands;
			track_o : out hex_char
		);
	end component node_52;
--sw  R1 ['68W02'] 
--dw  R1 [] 
--sc  R1 [] 
--lc  R1 [] 
	component route_0 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne1 : in hex_char;
			ne1_command : out routeCommands := RELEASE;
			s68W02_state : in hex_char;
			s68W02_command : out routeCommands := RELEASE;
			T02_state : in hex_char;
			T02_command : out routeCommands := RELEASE;
			C78_state : in hex_char;
			C78_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_0;
--sw  R2 ['68W02'] 
--dw  R2 [] 
--sc  R2 [] 
--lc  R2 [] 
	component route_1 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne7 : in hex_char;
			ne7_command : out routeCommands := RELEASE;
			s68W02_state : in hex_char;
			s68W02_command : out routeCommands := RELEASE;
			T06_state : in hex_char;
			T06_command : out routeCommands := RELEASE;
			J43_state : in hex_char;
			J43_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_1;
--sw  R3 ['69W04'] 
--dw  R3 [] 
--sc  R3 [] 
--lc  R3 [] 
	component route_2 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne14 : in hex_char;
			ne14_command : out routeCommands := RELEASE;
			track_ne52 : in hex_char;
			ne52_command : out routeCommands := RELEASE;
			s69W04_state : in hex_char;
			s69W04_command : out routeCommands := RELEASE;
			T08_state : in hex_char;
			T08_command : out routeCommands := RELEASE;
			S146_state : in hex_char;
			S146_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_2;
--sw  R4 ['71W02'] 
--dw  R4 [] 
--sc  R4 [] 
--lc  R4 [] 
	component route_3 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne47 : in hex_char;
			ne47_command : out routeCommands := RELEASE;
			track_ne48 : in hex_char;
			ne48_command : out routeCommands := RELEASE;
			s71W02_state : in hex_char;
			s71W02_command : out routeCommands := RELEASE;
			T12_state : in hex_char;
			T12_command : out routeCommands := RELEASE;
			L29_state : in hex_char;
			L29_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_3;
--sw  R5 ['Sw09', 'Sw04'] 
--dw  R5 ['Sw05'] 
--sc  R5 [] 
--lc  R5 [] 
	component route_4 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne84 : in hex_char;
			ne84_command : out routeCommands := RELEASE;
			track_ne82 : in hex_char;
			ne82_command : out routeCommands := RELEASE;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			T14_state : in hex_char;
			T14_command : out routeCommands := RELEASE;
			C100_state : in hex_char;
			C100_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_4;
--sw  R6 ['71W01', '71W02', 'Sw41'] 
--dw  R6 ['Sw05'] 
--sc  R6 [] 
--lc  R6 [] 
	component route_5 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne84 : in hex_char;
			ne84_command : out routeCommands := RELEASE;
			track_ne85 : in hex_char;
			ne85_command : out routeCommands := RELEASE;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			track_ne44 : in hex_char;
			ne44_command : out routeCommands := RELEASE;
			s71W01_state : in hex_char;
			s71W01_command : out routeCommands := RELEASE;
			s71W02_state : in hex_char;
			s71W02_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			T14_state : in hex_char;
			T14_command : out routeCommands := RELEASE;
			S105_state : in hex_char;
			S105_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_5;
--sw  R7 ['Sw08', 'Sw09', 'Sw12'] 
--dw  R7 [] 
--sc  R7 [] 
--lc  R7 [] 
	component route_6 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne89 : in hex_char;
			ne89_command : out routeCommands := RELEASE;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			T20_state : in hex_char;
			T20_command : out routeCommands := RELEASE;
			S97_state : in hex_char;
			S97_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_6;
--sw  R8 ['Sw08', 'Sw09', 'Sw12', 'Sw13'] 
--dw  R8 [] 
--sc  R8 [] 
--lc  R8 [] 
	component route_7 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne90 : in hex_char;
			ne90_command : out routeCommands := RELEASE;
			track_ne91 : in hex_char;
			ne91_command : out routeCommands := RELEASE;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			Sw13_state : in hex_char;
			Sw13_command : out routeCommands := RELEASE;
			T22_state : in hex_char;
			T22_command : out routeCommands := RELEASE;
			S97_state : in hex_char;
			S97_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_7;
--sw  R9 [] 
--dw  R9 [] 
--sc  R9 [] 
--lc  R9 [] 
	component route_8 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne105 : in hex_char;
			ne105_command : out routeCommands := RELEASE;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			track_ne96 : in hex_char;
			ne96_command : out routeCommands := RELEASE;
			T24_state : in hex_char;
			T24_command : out routeCommands := RELEASE;
			P70_state : in hex_char;
			P70_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_8;
--sw  R10 [] 
--dw  R10 [] 
--sc  R10 [] 
--lc  R10 [] 
	component route_9 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne4 : in hex_char;
			ne4_command : out routeCommands := RELEASE;
			track_ne106 : in hex_char;
			ne106_command : out routeCommands := RELEASE;
			L25_state : in hex_char;
			L25_command : out routeCommands := RELEASE;
			L42_state : in hex_char;
			L42_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_9;
--sw  R11 [] 
--dw  R11 [] 
--sc  R11 [] 
--lc  R11 [] 
	component route_10 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne26 : in hex_char;
			ne26_command : out routeCommands := RELEASE;
			track_ne65 : in hex_char;
			ne65_command : out routeCommands := RELEASE;
			L27_state : in hex_char;
			L27_command : out routeCommands := RELEASE;
			L30_state : in hex_char;
			L30_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_10;
--sw  R12 [] 
--dw  R12 [] 
--sc  R12 [] 
--lc  R12 [] 
	component route_11 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne44 : in hex_char;
			ne44_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			L28_state : in hex_char;
			L28_command : out routeCommands := RELEASE;
			L40_state : in hex_char;
			L40_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_11;
--sw  R13 ['71W01'] 
--dw  R13 [] 
--sc  R13 [] 
--lc  R13 [] 
	component route_12 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne65 : in hex_char;
			ne65_command : out routeCommands := RELEASE;
			track_ne102 : in hex_char;
			ne102_command : out routeCommands := RELEASE;
			s71W01_state : in hex_char;
			s71W01_command : out routeCommands := RELEASE;
			L30_state : in hex_char;
			L30_command : out routeCommands := RELEASE;
			C104_state : in hex_char;
			C104_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_12;
--sw  R14 ['Sw06'] 
--dw  R14 [] 
--sc  R14 ['Sw03'] 
--lc  R14 [] 
	component route_13 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne70 : in hex_char;
			ne70_command : out routeCommands := RELEASE;
			track_ne104 : in hex_char;
			ne104_command : out routeCommands := RELEASE;
			track_ne21 : in hex_char;
			ne21_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			L32_state : in hex_char;
			L32_command : out routeCommands := RELEASE;
			P73_state : in hex_char;
			P73_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_13;
--sw  R15 [] 
--dw  R15 [] 
--sc  R15 [] 
--lc  R15 [] 
	component route_14 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			track_ne93 : in hex_char;
			ne93_command : out routeCommands := RELEASE;
			L33_state : in hex_char;
			L33_command : out routeCommands := RELEASE;
			L34_state : in hex_char;
			L34_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_14;
--sw  R16 [] 
--dw  R16 [] 
--sc  R16 [] 
--lc  R16 [] 
	component route_15 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne93 : in hex_char;
			ne93_command : out routeCommands := RELEASE;
			track_ne96 : in hex_char;
			ne96_command : out routeCommands := RELEASE;
			L34_state : in hex_char;
			L34_command : out routeCommands := RELEASE;
			P71_state : in hex_char;
			P71_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_15;
--sw  R17 [] 
--dw  R17 [] 
--sc  R17 [] 
--lc  R17 [] 
	component route_16 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne95 : in hex_char;
			ne95_command : out routeCommands := RELEASE;
			L35_state : in hex_char;
			L35_command : out routeCommands := RELEASE;
			X50_state : in hex_char;
			X50_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_16;
--sw  R18 [] 
--dw  R18 [] 
--sc  R18 [] 
--lc  R18 [] 
	component route_17 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne97 : in hex_char;
			ne97_command : out routeCommands := RELEASE;
			track_ne94 : in hex_char;
			ne94_command : out routeCommands := RELEASE;
			L37_state : in hex_char;
			L37_command : out routeCommands := RELEASE;
			S135_state : in hex_char;
			S135_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_17;
--sw  R19 [] 
--dw  R19 [] 
--sc  R19 [] 
--lc  R19 [] 
	component route_18 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			track_ne105 : in hex_char;
			ne105_command : out routeCommands := RELEASE;
			L38_state : in hex_char;
			L38_command : out routeCommands := RELEASE;
			T23_state : in hex_char;
			T23_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_18;
--sw  R20 ['Sw41'] 
--dw  R20 [] 
--sc  R20 [] 
--lc  R20 [] 
	component route_19 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			L40_state : in hex_char;
			L40_command : out routeCommands := RELEASE;
			S139_state : in hex_char;
			S139_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_19;
--sw  R21 ['70W01'] 
--dw  R21 [] 
--sc  R21 [] 
--lc  R21 [] 
	component route_20 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne103 : in hex_char;
			ne103_command : out routeCommands := RELEASE;
			track_ne64 : in hex_char;
			ne64_command : out routeCommands := RELEASE;
			s70W01_state : in hex_char;
			s70W01_command : out routeCommands := RELEASE;
			L41_state : in hex_char;
			L41_command : out routeCommands := RELEASE;
			S90_state : in hex_char;
			S90_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_20;
--sw  R22 [] 
--dw  R22 [] 
--sc  R22 [] 
--lc  R22 [] 
	component route_21 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne106 : in hex_char;
			ne106_command : out routeCommands := RELEASE;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			L42_state : in hex_char;
			L42_command : out routeCommands := RELEASE;
			P68_state : in hex_char;
			P68_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_21;
--sw  R23 ['68W02'] 
--dw  R23 [] 
--sc  R23 [] 
--lc  R23 [] 
	component route_22 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne7 : in hex_char;
			ne7_command : out routeCommands := RELEASE;
			track_ne9 : in hex_char;
			ne9_command : out routeCommands := RELEASE;
			s68W02_state : in hex_char;
			s68W02_command : out routeCommands := RELEASE;
			J43_state : in hex_char;
			J43_command : out routeCommands := RELEASE;
			J46_state : in hex_char;
			J46_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_22;
--sw  R24 [] 
--dw  R24 [] 
--sc  R24 [] 
--lc  R24 [] 
	component route_23 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne9 : in hex_char;
			ne9_command : out routeCommands := RELEASE;
			track_ne95 : in hex_char;
			ne95_command : out routeCommands := RELEASE;
			J46_state : in hex_char;
			J46_command : out routeCommands := RELEASE;
			L35_state : in hex_char;
			L35_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_23;
--sw  R25 ['69W03', '69W04'] 
--dw  R25 [] 
--sc  R25 [] 
--lc  R25 ['Lc01'] 
	component route_24 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne95 : in hex_char;
			ne95_command : out routeCommands := RELEASE;
			track_ne59 : in hex_char;
			ne59_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			s69W03_state : in hex_char;
			s69W03_command : out routeCommands := RELEASE;
			s69W04_state : in hex_char;
			s69W04_command : out routeCommands := RELEASE;
			X50_state : in hex_char;
			X50_command : out routeCommands := RELEASE;
			S83_state : in hex_char;
			S83_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_24;
--sw  R26 ['68W02'] 
--dw  R26 [] 
--sc  R26 [] 
--lc  R26 ['Lc01'] 
	component route_25 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne95 : in hex_char;
			ne95_command : out routeCommands := RELEASE;
			track_ne9 : in hex_char;
			ne9_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			s68W02_state : in hex_char;
			s68W02_command : out routeCommands := RELEASE;
			X51_state : in hex_char;
			X51_command : out routeCommands := RELEASE;
			S80_state : in hex_char;
			S80_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_25;
--sw  R27 ['70W02'] 
--dw  R27 [] 
--sc  R27 [] 
--lc  R27 [] 
	component route_26 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne23 : in hex_char;
			ne23_command : out routeCommands := RELEASE;
			track_ne26 : in hex_char;
			ne26_command : out routeCommands := RELEASE;
			s70W02_state : in hex_char;
			s70W02_command : out routeCommands := RELEASE;
			P60_state : in hex_char;
			P60_command : out routeCommands := RELEASE;
			L27_state : in hex_char;
			L27_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_26;
--sw  R28 [] 
--dw  R28 [] 
--sc  R28 [] 
--lc  R28 [] 
	component route_27 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne24 : in hex_char;
			ne24_command : out routeCommands := RELEASE;
			track_ne64 : in hex_char;
			ne64_command : out routeCommands := RELEASE;
			track_ne103 : in hex_char;
			ne103_command : out routeCommands := RELEASE;
			track_ne67 : in hex_char;
			ne67_command : out routeCommands := RELEASE;
			P63_state : in hex_char;
			P63_command : out routeCommands := RELEASE;
			P64_state : in hex_char;
			P64_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_27;
--sw  R29 [] 
--dw  R29 [] 
--sc  R29 [] 
--lc  R29 [] 
	component route_28 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne67 : in hex_char;
			ne67_command : out routeCommands := RELEASE;
			track_ne70 : in hex_char;
			ne70_command : out routeCommands := RELEASE;
			P64_state : in hex_char;
			P64_command : out routeCommands := RELEASE;
			L32_state : in hex_char;
			L32_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_28;
--sw  R30 [] 
--dw  R30 [] 
--sc  R30 [] 
--lc  R30 [] 
	component route_29 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne67 : in hex_char;
			ne67_command : out routeCommands := RELEASE;
			track_ne103 : in hex_char;
			ne103_command : out routeCommands := RELEASE;
			P65_state : in hex_char;
			P65_command : out routeCommands := RELEASE;
			L41_state : in hex_char;
			L41_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_29;
--sw  R31 [] 
--dw  R31 [] 
--sc  R31 [] 
--lc  R31 [] 
	component route_30 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			track_ne97 : in hex_char;
			ne97_command : out routeCommands := RELEASE;
			P68_state : in hex_char;
			P68_command : out routeCommands := RELEASE;
			L37_state : in hex_char;
			L37_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_30;
--sw  R32 [] 
--dw  R32 [] 
--sc  R32 [] 
--lc  R32 [] 
	component route_31 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			track_ne106 : in hex_char;
			ne106_command : out routeCommands := RELEASE;
			track_ne4 : in hex_char;
			ne4_command : out routeCommands := RELEASE;
			P69_state : in hex_char;
			P69_command : out routeCommands := RELEASE;
			T03_state : in hex_char;
			T03_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_31;
--sw  R33 ['Sw06'] 
--dw  R33 [] 
--sc  R33 [] 
--lc  R33 [] 
	component route_32 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne96 : in hex_char;
			ne96_command : out routeCommands := RELEASE;
			track_ne93 : in hex_char;
			ne93_command : out routeCommands := RELEASE;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			P70_state : in hex_char;
			P70_command : out routeCommands := RELEASE;
			S110_state : in hex_char;
			S110_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_32;
--sw  R34 [] 
--dw  R34 [] 
--sc  R34 [] 
--lc  R34 [] 
	component route_33 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne96 : in hex_char;
			ne96_command : out routeCommands := RELEASE;
			track_ne98 : in hex_char;
			ne98_command : out routeCommands := RELEASE;
			P71_state : in hex_char;
			P71_command : out routeCommands := RELEASE;
			L38_state : in hex_char;
			L38_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_33;
--sw  R35 [] 
--dw  R35 [] 
--sc  R35 [] 
--lc  R35 [] 
	component route_34 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne21 : in hex_char;
			ne21_command : out routeCommands := RELEASE;
			P72_state : in hex_char;
			P72_command : out routeCommands := RELEASE;
			S144_state : in hex_char;
			S144_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_34;
--sw  R36 ['Sw06'] 
--dw  R36 ['Sw07'] 
--sc  R36 [] 
--lc  R36 [] 
	component route_35 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne21 : in hex_char;
			ne21_command : out routeCommands := RELEASE;
			track_ne79 : in hex_char;
			ne79_command : out routeCommands := RELEASE;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			P73_state : in hex_char;
			P73_command : out routeCommands := RELEASE;
			L33_state : in hex_char;
			L33_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_35;
--sw  R37 [] 
--dw  R37 ['Sw07'] 
--sc  R37 [] 
--lc  R37 [] 
	component route_36 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne21 : in hex_char;
			ne21_command : out routeCommands := RELEASE;
			track_ne94 : in hex_char;
			ne94_command : out routeCommands := RELEASE;
			track_ne97 : in hex_char;
			ne97_command : out routeCommands := RELEASE;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			P73_state : in hex_char;
			P73_command : out routeCommands := RELEASE;
			P69_state : in hex_char;
			P69_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_36;
--sw  R38 ['68W02'] 
--dw  R38 [] 
--sc  R38 [] 
--lc  R38 [] 
	component route_37 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne1 : in hex_char;
			ne1_command : out routeCommands := RELEASE;
			track_ne9 : in hex_char;
			ne9_command : out routeCommands := RELEASE;
			s68W02_state : in hex_char;
			s68W02_command : out routeCommands := RELEASE;
			C78_state : in hex_char;
			C78_command : out routeCommands := RELEASE;
			J46_state : in hex_char;
			J46_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_37;
--sw  R39 ['68W02'] 
--dw  R39 [] 
--sc  R39 [] 
--lc  R39 [] 
	component route_38 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne9 : in hex_char;
			ne9_command : out routeCommands := RELEASE;
			track_ne1 : in hex_char;
			ne1_command : out routeCommands := RELEASE;
			s68W02_state : in hex_char;
			s68W02_command : out routeCommands := RELEASE;
			S80_state : in hex_char;
			S80_command : out routeCommands := RELEASE;
			T01_state : in hex_char;
			T01_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_38;
--sw  R40 ['68W02'] 
--dw  R40 [] 
--sc  R40 [] 
--lc  R40 [] 
	component route_39 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne9 : in hex_char;
			ne9_command : out routeCommands := RELEASE;
			track_ne7 : in hex_char;
			ne7_command : out routeCommands := RELEASE;
			s68W02_state : in hex_char;
			s68W02_command : out routeCommands := RELEASE;
			S80_state : in hex_char;
			S80_command : out routeCommands := RELEASE;
			T05_state : in hex_char;
			T05_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_39;
--sw  R41 ['69W03'] 
--dw  R41 [] 
--sc  R41 [] 
--lc  R41 ['Lc01'] 
	component route_40 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne17 : in hex_char;
			ne17_command : out routeCommands := RELEASE;
			track_ne59 : in hex_char;
			ne59_command : out routeCommands := RELEASE;
			track_ne95 : in hex_char;
			ne95_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			s69W03_state : in hex_char;
			s69W03_command : out routeCommands := RELEASE;
			C82_state : in hex_char;
			C82_command : out routeCommands := RELEASE;
			X51_state : in hex_char;
			X51_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_40;
--sw  R42 ['69W03', '69W04'] 
--dw  R42 [] 
--sc  R42 [] 
--lc  R42 [] 
	component route_41 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne59 : in hex_char;
			ne59_command : out routeCommands := RELEASE;
			track_ne11 : in hex_char;
			ne11_command : out routeCommands := RELEASE;
			track_ne52 : in hex_char;
			ne52_command : out routeCommands := RELEASE;
			s69W03_state : in hex_char;
			s69W03_command : out routeCommands := RELEASE;
			s69W04_state : in hex_char;
			s69W04_command : out routeCommands := RELEASE;
			S83_state : in hex_char;
			S83_command : out routeCommands := RELEASE;
			S146_state : in hex_char;
			S146_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_41;
--sw  R43 ['69W03', 'Sw06'] 
--dw  R43 [] 
--sc  R43 [] 
--lc  R43 [] 
	component route_42 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne59 : in hex_char;
			ne59_command : out routeCommands := RELEASE;
			track_ne17 : in hex_char;
			ne17_command : out routeCommands := RELEASE;
			s69W03_state : in hex_char;
			s69W03_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			S83_state : in hex_char;
			S83_command : out routeCommands := RELEASE;
			C109_state : in hex_char;
			C109_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_42;
--sw  R44 ['69W03', '69W04'] 
--dw  R44 [] 
--sc  R44 [] 
--lc  R44 ['Lc01'] 
	component route_43 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne52 : in hex_char;
			ne52_command : out routeCommands := RELEASE;
			track_ne11 : in hex_char;
			ne11_command : out routeCommands := RELEASE;
			track_ne59 : in hex_char;
			ne59_command : out routeCommands := RELEASE;
			track_ne95 : in hex_char;
			ne95_command : out routeCommands := RELEASE;
			Lc01_state : in hex_char;
			Lc01_command : out routeCommands := RELEASE;
			s69W03_state : in hex_char;
			s69W03_command : out routeCommands := RELEASE;
			s69W04_state : in hex_char;
			s69W04_command : out routeCommands := RELEASE;
			S86_state : in hex_char;
			S86_command : out routeCommands := RELEASE;
			X51_state : in hex_char;
			X51_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_43;
--sw  R45 ['69W04'] 
--dw  R45 [] 
--sc  R45 [] 
--lc  R45 [] 
	component route_44 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne52 : in hex_char;
			ne52_command : out routeCommands := RELEASE;
			track_ne14 : in hex_char;
			ne14_command : out routeCommands := RELEASE;
			s69W04_state : in hex_char;
			s69W04_command : out routeCommands := RELEASE;
			S86_state : in hex_char;
			S86_command : out routeCommands := RELEASE;
			T07_state : in hex_char;
			T07_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_44;
--sw  R46 [] 
--dw  R46 [] 
--sc  R46 [] 
--lc  R46 [] 
	component route_45 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne23 : in hex_char;
			ne23_command : out routeCommands := RELEASE;
			track_ne64 : in hex_char;
			ne64_command : out routeCommands := RELEASE;
			track_ne103 : in hex_char;
			ne103_command : out routeCommands := RELEASE;
			track_ne67 : in hex_char;
			ne67_command : out routeCommands := RELEASE;
			B89_state : in hex_char;
			B89_command : out routeCommands := RELEASE;
			P64_state : in hex_char;
			P64_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_45;
--sw  R47 ['70W01', '70W02'] 
--dw  R47 [] 
--sc  R47 [] 
--lc  R47 [] 
	component route_46 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne64 : in hex_char;
			ne64_command : out routeCommands := RELEASE;
			track_ne23 : in hex_char;
			ne23_command : out routeCommands := RELEASE;
			s70W01_state : in hex_char;
			s70W01_command : out routeCommands := RELEASE;
			s70W02_state : in hex_char;
			s70W02_command : out routeCommands := RELEASE;
			S90_state : in hex_char;
			S90_command : out routeCommands := RELEASE;
			P60_state : in hex_char;
			P60_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_46;
--sw  R48 ['70W01', '70W02'] 
--dw  R48 [] 
--sc  R48 [] 
--lc  R48 [] 
	component route_47 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne64 : in hex_char;
			ne64_command : out routeCommands := RELEASE;
			track_ne24 : in hex_char;
			ne24_command : out routeCommands := RELEASE;
			s70W01_state : in hex_char;
			s70W01_command : out routeCommands := RELEASE;
			s70W02_state : in hex_char;
			s70W02_command : out routeCommands := RELEASE;
			S90_state : in hex_char;
			S90_command : out routeCommands := RELEASE;
			B92_state : in hex_char;
			B92_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_47;
--sw  R49 ['70W02'] 
--dw  R49 [] 
--sc  R49 [] 
--lc  R49 [] 
	component route_48 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne24 : in hex_char;
			ne24_command : out routeCommands := RELEASE;
			track_ne26 : in hex_char;
			ne26_command : out routeCommands := RELEASE;
			s70W02_state : in hex_char;
			s70W02_command : out routeCommands := RELEASE;
			B92_state : in hex_char;
			B92_command : out routeCommands := RELEASE;
			L27_state : in hex_char;
			L27_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_48;
--sw  R50 ['70W02'] 
--dw  R50 [] 
--sc  R50 [] 
--lc  R50 [] 
	component route_49 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne26 : in hex_char;
			ne26_command : out routeCommands := RELEASE;
			track_ne23 : in hex_char;
			ne23_command : out routeCommands := RELEASE;
			s70W02_state : in hex_char;
			s70W02_command : out routeCommands := RELEASE;
			S93_state : in hex_char;
			S93_command : out routeCommands := RELEASE;
			B89_state : in hex_char;
			B89_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_49;
--sw  R51 ['70W02'] 
--dw  R51 [] 
--sc  R51 [] 
--lc  R51 [] 
	component route_50 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne26 : in hex_char;
			ne26_command : out routeCommands := RELEASE;
			track_ne24 : in hex_char;
			ne24_command : out routeCommands := RELEASE;
			s70W02_state : in hex_char;
			s70W02_command : out routeCommands := RELEASE;
			S93_state : in hex_char;
			S93_command : out routeCommands := RELEASE;
			P63_state : in hex_char;
			P63_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_50;
--sw  R52 ['Sw08', 'Sw12'] 
--dw  R52 [] 
--sc  R52 [] 
--lc  R52 [] 
	component route_51 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne83 : in hex_char;
			ne83_command : out routeCommands := RELEASE;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			C95_state : in hex_char;
			C95_command : out routeCommands := RELEASE;
			S122_state : in hex_char;
			S122_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_51;
--sw  R53 ['Sw08', 'Sw12'] 
--dw  R53 [] 
--sc  R53 [] 
--lc  R53 [] 
	component route_52 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne29 : in hex_char;
			ne29_command : out routeCommands := RELEASE;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			B96_state : in hex_char;
			B96_command : out routeCommands := RELEASE;
			S122_state : in hex_char;
			S122_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_52;
--sw  R54 ['Sw08', 'Sw09', 'Sw41'] 
--dw  R54 [] 
--sc  R54 [] 
--lc  R54 [] 
	component route_53 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			track_ne29 : in hex_char;
			ne29_command : out routeCommands := RELEASE;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			S97_state : in hex_char;
			S97_command : out routeCommands := RELEASE;
			C138_state : in hex_char;
			C138_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_53;
--sw  R55 ['Sw08', 'Sw04'] 
--dw  R55 [] 
--sc  R55 [] 
--lc  R55 [] 
	component route_54 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			track_ne83 : in hex_char;
			ne83_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			S97_state : in hex_char;
			S97_command : out routeCommands := RELEASE;
			C114_state : in hex_char;
			C114_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_54;
--sw  R56 ['Sw09', 'Sw41'] 
--dw  R56 [] 
--sc  R56 [] 
--lc  R56 [] 
	component route_55 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			C100_state : in hex_char;
			C100_command : out routeCommands := RELEASE;
			C138_state : in hex_char;
			C138_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_55;
--sw  R57 ['Sw08'] 
--dw  R57 [] 
--sc  R57 [] 
--lc  R57 [] 
	component route_56 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne29 : in hex_char;
			ne29_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			B101_state : in hex_char;
			B101_command : out routeCommands := RELEASE;
			B96_state : in hex_char;
			B96_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_56;
--sw  R58 ['Sw09', 'Sw04'] 
--dw  R58 [] 
--sc  R58 [] 
--lc  R58 [] 
	component route_57 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			S102_state : in hex_char;
			S102_command : out routeCommands := RELEASE;
			S115_state : in hex_char;
			S115_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_57;
--sw  R59 ['Sw09'] 
--dw  R59 [] 
--sc  R59 [] 
--lc  R59 [] 
	component route_58 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			track_ne29 : in hex_char;
			ne29_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			S102_state : in hex_char;
			S102_command : out routeCommands := RELEASE;
			B101_state : in hex_char;
			B101_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_58;
--sw  R60 ['71W01'] 
--dw  R60 [] 
--sc  R60 [] 
--lc  R60 [] 
	component route_59 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne102 : in hex_char;
			ne102_command : out routeCommands := RELEASE;
			track_ne44 : in hex_char;
			ne44_command : out routeCommands := RELEASE;
			s71W01_state : in hex_char;
			s71W01_command : out routeCommands := RELEASE;
			C104_state : in hex_char;
			C104_command : out routeCommands := RELEASE;
			L28_state : in hex_char;
			L28_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_59;
--sw  R61 ['71W01', '71W02'] 
--dw  R61 [] 
--sc  R61 [] 
--lc  R61 [] 
	component route_60 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne44 : in hex_char;
			ne44_command : out routeCommands := RELEASE;
			track_ne43 : in hex_char;
			ne43_command : out routeCommands := RELEASE;
			track_ne48 : in hex_char;
			ne48_command : out routeCommands := RELEASE;
			s71W01_state : in hex_char;
			s71W01_command : out routeCommands := RELEASE;
			s71W02_state : in hex_char;
			s71W02_command : out routeCommands := RELEASE;
			S105_state : in hex_char;
			S105_command : out routeCommands := RELEASE;
			L29_state : in hex_char;
			L29_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_60;
--sw  R62 ['70W02', '71W01'] 
--dw  R62 [] 
--sc  R62 [] 
--lc  R62 [] 
	component route_61 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne44 : in hex_char;
			ne44_command : out routeCommands := RELEASE;
			track_ne102 : in hex_char;
			ne102_command : out routeCommands := RELEASE;
			track_ne65 : in hex_char;
			ne65_command : out routeCommands := RELEASE;
			track_ne26 : in hex_char;
			ne26_command : out routeCommands := RELEASE;
			s70W02_state : in hex_char;
			s70W02_command : out routeCommands := RELEASE;
			s71W01_state : in hex_char;
			s71W01_command : out routeCommands := RELEASE;
			S105_state : in hex_char;
			S105_command : out routeCommands := RELEASE;
			S93_state : in hex_char;
			S93_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_61;
--sw  R63 ['Sw06'] 
--dw  R63 [] 
--sc  R63 [] 
--lc  R63 [] 
	component route_62 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne17 : in hex_char;
			ne17_command : out routeCommands := RELEASE;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			C109_state : in hex_char;
			C109_command : out routeCommands := RELEASE;
			L33_state : in hex_char;
			L33_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_62;
--sw  R64 ['69W03', 'Sw06'] 
--dw  R64 [] 
--sc  R64 [] 
--lc  R64 [] 
	component route_63 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			track_ne17 : in hex_char;
			ne17_command : out routeCommands := RELEASE;
			s69W03_state : in hex_char;
			s69W03_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			S110_state : in hex_char;
			S110_command : out routeCommands := RELEASE;
			C82_state : in hex_char;
			C82_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_63;
--sw  R65 ['Sw06'] 
--dw  R65 ['Sw07'] 
--sc  R65 [] 
--lc  R65 [] 
	component route_64 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			track_ne79 : in hex_char;
			ne79_command : out routeCommands := RELEASE;
			track_ne77 : in hex_char;
			ne77_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			S110_state : in hex_char;
			S110_command : out routeCommands := RELEASE;
			B133_state : in hex_char;
			B133_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_64;
--sw  R66 ['Sw06'] 
--dw  R66 ['Sw07'] 
--sc  R66 [] 
--lc  R66 [] 
	component route_65 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			track_ne79 : in hex_char;
			ne79_command : out routeCommands := RELEASE;
			track_ne21 : in hex_char;
			ne21_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			S110_state : in hex_char;
			S110_command : out routeCommands := RELEASE;
			P72_state : in hex_char;
			P72_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_65;
--sw  R67 ['Sw09', 'Sw04'] 
--dw  R67 [] 
--sc  R67 [] 
--lc  R67 [] 
	component route_66 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne83 : in hex_char;
			ne83_command : out routeCommands := RELEASE;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			C114_state : in hex_char;
			C114_command : out routeCommands := RELEASE;
			C100_state : in hex_char;
			C100_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_66;
--sw  R68 ['Sw08', 'Sw04'] 
--dw  R68 [] 
--sc  R68 [] 
--lc  R68 [] 
	component route_67 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			track_ne83 : in hex_char;
			ne83_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			S115_state : in hex_char;
			S115_command : out routeCommands := RELEASE;
			C95_state : in hex_char;
			C95_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_67;
--sw  R69 ['Sw04'] 
--dw  R69 ['Sw05'] 
--sc  R69 [] 
--lc  R69 [] 
	component route_68 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			track_ne82 : in hex_char;
			ne82_command : out routeCommands := RELEASE;
			track_ne41 : in hex_char;
			ne41_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			S115_state : in hex_char;
			S115_command : out routeCommands := RELEASE;
			P58_state : in hex_char;
			P58_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_68;
--sw  R70 ['Sw04'] 
--dw  R70 ['Sw05'] 
--sc  R70 [] 
--lc  R70 [] 
	component route_69 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			track_ne82 : in hex_char;
			ne82_command : out routeCommands := RELEASE;
			track_ne84 : in hex_char;
			ne84_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			S115_state : in hex_char;
			S115_command : out routeCommands := RELEASE;
			T13_state : in hex_char;
			T13_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_69;
--sw  R71 ['Sw11'] 
--dw  R71 [] 
--sc  R71 [] 
--lc  R71 [] 
	component route_70 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne88 : in hex_char;
			ne88_command : out routeCommands := RELEASE;
			track_ne86 : in hex_char;
			ne86_command : out routeCommands := RELEASE;
			Sw11_state : in hex_char;
			Sw11_command : out routeCommands := RELEASE;
			C118_state : in hex_char;
			C118_command : out routeCommands := RELEASE;
			T15_state : in hex_char;
			T15_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_70;
--sw  R72 ['Sw11'] 
--dw  R72 [] 
--sc  R72 [] 
--lc  R72 [] 
	component route_71 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne86 : in hex_char;
			ne86_command : out routeCommands := RELEASE;
			track_ne88 : in hex_char;
			ne88_command : out routeCommands := RELEASE;
			Sw11_state : in hex_char;
			Sw11_command : out routeCommands := RELEASE;
			S119_state : in hex_char;
			S119_command : out routeCommands := RELEASE;
			T17_state : in hex_char;
			T17_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_71;
--sw  R73 ['Sw08', 'Sw09', 'Sw12', 'Sw11', 'Sw13'] 
--dw  R73 [] 
--sc  R73 [] 
--lc  R73 [] 
	component route_72 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne86 : in hex_char;
			ne86_command : out routeCommands := RELEASE;
			track_ne87 : in hex_char;
			ne87_command : out routeCommands := RELEASE;
			track_ne91 : in hex_char;
			ne91_command : out routeCommands := RELEASE;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			Sw08_state : in hex_char;
			Sw08_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			Sw11_state : in hex_char;
			Sw11_command : out routeCommands := RELEASE;
			Sw13_state : in hex_char;
			Sw13_command : out routeCommands := RELEASE;
			S119_state : in hex_char;
			S119_command : out routeCommands := RELEASE;
			S97_state : in hex_char;
			S97_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_72;
--sw  R74 ['Sw12'] 
--dw  R74 [] 
--sc  R74 [] 
--lc  R74 [] 
	component route_73 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			track_ne89 : in hex_char;
			ne89_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			S122_state : in hex_char;
			S122_command : out routeCommands := RELEASE;
			T19_state : in hex_char;
			T19_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_73;
--sw  R75 ['Sw12', 'Sw11', 'Sw13'] 
--dw  R75 [] 
--sc  R75 [] 
--lc  R75 [] 
	component route_74 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			track_ne91 : in hex_char;
			ne91_command : out routeCommands := RELEASE;
			track_ne87 : in hex_char;
			ne87_command : out routeCommands := RELEASE;
			track_ne86 : in hex_char;
			ne86_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			Sw11_state : in hex_char;
			Sw11_command : out routeCommands := RELEASE;
			Sw13_state : in hex_char;
			Sw13_command : out routeCommands := RELEASE;
			S122_state : in hex_char;
			S122_command : out routeCommands := RELEASE;
			T15_state : in hex_char;
			T15_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_74;
--sw  R76 ['Sw12', 'Sw13'] 
--dw  R76 [] 
--sc  R76 [] 
--lc  R76 [] 
	component route_75 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne30 : in hex_char;
			ne30_command : out routeCommands := RELEASE;
			track_ne91 : in hex_char;
			ne91_command : out routeCommands := RELEASE;
			track_ne90 : in hex_char;
			ne90_command : out routeCommands := RELEASE;
			Sw12_state : in hex_char;
			Sw12_command : out routeCommands := RELEASE;
			Sw13_state : in hex_char;
			Sw13_command : out routeCommands := RELEASE;
			S122_state : in hex_char;
			S122_command : out routeCommands := RELEASE;
			T21_state : in hex_char;
			T21_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_75;
--sw  R77 ['Sw09', 'Sw04'] 
--dw  R77 ['Sw05'] 
--sc  R77 [] 
--lc  R77 [] 
	component route_76 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne41 : in hex_char;
			ne41_command : out routeCommands := RELEASE;
			track_ne82 : in hex_char;
			ne82_command : out routeCommands := RELEASE;
			track_ne32 : in hex_char;
			ne32_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw04_state : in hex_char;
			Sw04_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			B130_state : in hex_char;
			B130_command : out routeCommands := RELEASE;
			C100_state : in hex_char;
			C100_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_76;
--sw  R78 ['71W01', '71W02', 'Sw41'] 
--dw  R78 ['Sw05'] 
--sc  R78 [] 
--lc  R78 [] 
	component route_77 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne41 : in hex_char;
			ne41_command : out routeCommands := RELEASE;
			track_ne85 : in hex_char;
			ne85_command : out routeCommands := RELEASE;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			track_ne44 : in hex_char;
			ne44_command : out routeCommands := RELEASE;
			s71W01_state : in hex_char;
			s71W01_command : out routeCommands := RELEASE;
			s71W02_state : in hex_char;
			s71W02_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			B130_state : in hex_char;
			B130_command : out routeCommands := RELEASE;
			S105_state : in hex_char;
			S105_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_77;
--sw  R79 [] 
--dw  R79 ['Sw05'] 
--sc  R79 [] 
--lc  R79 [] 
	component route_78 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne85 : in hex_char;
			ne85_command : out routeCommands := RELEASE;
			track_ne41 : in hex_char;
			ne41_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			S131_state : in hex_char;
			S131_command : out routeCommands := RELEASE;
			P58_state : in hex_char;
			P58_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_78;
--sw  R80 [] 
--dw  R80 ['Sw05'] 
--sc  R80 [] 
--lc  R80 [] 
	component route_79 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne85 : in hex_char;
			ne85_command : out routeCommands := RELEASE;
			track_ne84 : in hex_char;
			ne84_command : out routeCommands := RELEASE;
			Sw05_state : in hex_char;
			Sw05_command : out routeCommands := RELEASE;
			S131_state : in hex_char;
			S131_command : out routeCommands := RELEASE;
			T13_state : in hex_char;
			T13_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_79;
--sw  R81 ['69W03', '69W04'] 
--dw  R81 [] 
--sc  R81 ['Sw03'] 
--lc  R81 [] 
	component route_80 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne77 : in hex_char;
			ne77_command : out routeCommands := RELEASE;
			track_ne52 : in hex_char;
			ne52_command : out routeCommands := RELEASE;
			s69W03_state : in hex_char;
			s69W03_command : out routeCommands := RELEASE;
			s69W04_state : in hex_char;
			s69W04_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			B133_state : in hex_char;
			B133_command : out routeCommands := RELEASE;
			S86_state : in hex_char;
			S86_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_80;
--sw  R82 [] 
--dw  R82 ['Sw07'] 
--sc  R82 [] 
--lc  R82 [] 
	component route_81 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne94 : in hex_char;
			ne94_command : out routeCommands := RELEASE;
			track_ne77 : in hex_char;
			ne77_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			S135_state : in hex_char;
			S135_command : out routeCommands := RELEASE;
			B133_state : in hex_char;
			B133_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_81;
--sw  R83 [] 
--dw  R83 ['Sw07'] 
--sc  R83 [] 
--lc  R83 [] 
	component route_82 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne94 : in hex_char;
			ne94_command : out routeCommands := RELEASE;
			track_ne21 : in hex_char;
			ne21_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			S135_state : in hex_char;
			S135_command : out routeCommands := RELEASE;
			P72_state : in hex_char;
			P72_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_82;
--sw  R84 ['71W01', '71W02', 'Sw41'] 
--dw  R84 [] 
--sc  R84 [] 
--lc  R84 [] 
	component route_83 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			track_ne101 : in hex_char;
			ne101_command : out routeCommands := RELEASE;
			track_ne44 : in hex_char;
			ne44_command : out routeCommands := RELEASE;
			s71W01_state : in hex_char;
			s71W01_command : out routeCommands := RELEASE;
			s71W02_state : in hex_char;
			s71W02_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			C138_state : in hex_char;
			C138_command : out routeCommands := RELEASE;
			S105_state : in hex_char;
			S105_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_83;
--sw  R85 ['Sw09', 'Sw41'] 
--dw  R85 [] 
--sc  R85 [] 
--lc  R85 [] 
	component route_84 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			track_ne110 : in hex_char;
			ne110_command : out routeCommands := RELEASE;
			Sw09_state : in hex_char;
			Sw09_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			S139_state : in hex_char;
			S139_command : out routeCommands := RELEASE;
			S102_state : in hex_char;
			S102_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_84;
--sw  R86 ['Sw41'] 
--dw  R86 [] 
--sc  R86 [] 
--lc  R86 [] 
	component route_85 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne100 : in hex_char;
			ne100_command : out routeCommands := RELEASE;
			track_ne85 : in hex_char;
			ne85_command : out routeCommands := RELEASE;
			Sw41_state : in hex_char;
			Sw41_command : out routeCommands := RELEASE;
			S139_state : in hex_char;
			S139_command : out routeCommands := RELEASE;
			S131_state : in hex_char;
			S131_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_85;
--sw  R87 [] 
--dw  R87 [] 
--sc  R87 [] 
--lc  R87 [] 
	component route_86 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne104 : in hex_char;
			ne104_command : out routeCommands := RELEASE;
			track_ne70 : in hex_char;
			ne70_command : out routeCommands := RELEASE;
			B143_state : in hex_char;
			B143_command : out routeCommands := RELEASE;
			L32_state : in hex_char;
			L32_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_86;
--sw  R88 [] 
--dw  R88 [] 
--sc  R88 ['Sw03'] 
--lc  R88 [] 
	component route_87 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne21 : in hex_char;
			ne21_command : out routeCommands := RELEASE;
			track_ne104 : in hex_char;
			ne104_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			S144_state : in hex_char;
			S144_command : out routeCommands := RELEASE;
			B143_state : in hex_char;
			B143_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_87;
--sw  R89 ['Sw06'] 
--dw  R89 ['Sw07'] 
--sc  R89 [] 
--lc  R89 [] 
	component route_88 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne77 : in hex_char;
			ne77_command : out routeCommands := RELEASE;
			track_ne79 : in hex_char;
			ne79_command : out routeCommands := RELEASE;
			track_ne78 : in hex_char;
			ne78_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			B145_state : in hex_char;
			B145_command : out routeCommands := RELEASE;
			L33_state : in hex_char;
			L33_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_88;
--sw  R90 [] 
--dw  R90 ['Sw07'] 
--sc  R90 [] 
--lc  R90 [] 
	component route_89 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne77 : in hex_char;
			ne77_command : out routeCommands := RELEASE;
			track_ne94 : in hex_char;
			ne94_command : out routeCommands := RELEASE;
			track_ne97 : in hex_char;
			ne97_command : out routeCommands := RELEASE;
			track_ne99 : in hex_char;
			ne99_command : out routeCommands := RELEASE;
			Sw07_state : in hex_char;
			Sw07_command : out routeCommands := RELEASE;
			B145_state : in hex_char;
			B145_command : out routeCommands := RELEASE;
			P69_state : in hex_char;
			P69_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_89;
--sw  R91 ['Sw06'] 
--dw  R91 [] 
--sc  R91 ['Sw03'] 
--lc  R91 [] 
	component route_90 is
		port(
			clock : in std_logic := '0';
			reset : in std_logic := '0';
			routeRequest : in hex_char;
			track_ne52 : in hex_char;
			ne52_command : out routeCommands := RELEASE;
			track_ne77 : in hex_char;
			ne77_command : out routeCommands := RELEASE;
			Sw06_state : in hex_char;
			Sw06_command : out routeCommands := RELEASE;
			Sw03_state : in hex_char;
			Sw03_command : out routeCommands := RELEASE;
			S146_state : in hex_char;
			S146_command : out routeCommands := RELEASE;
			B145_state : in hex_char;
			B145_command : out routeCommands := RELEASE;
			routeExecute : out hex_char
		);
	end component route_90;
	signal state_Lc01 : hex_char;
	signal state_68W02 , state_69W03 , state_69W04 , state_Sw06 , state_70W01 , state_70W02 , state_Sw08 , state_Sw09 , state_Sw12 , state_Sw04 , state_71W01 , state_71W02 , state_Sw11 , state_Sw13 , state_Sw41 : hex_char;
	signal state_Sw03 : hex_char;
	signal state_Sw05 , state_Sw07 : hex_char;
	signal state_T01 , state_T02 , state_C78 , state_T03 , state_L25 , state_T05 , state_T06 , state_J43 , state_J46 , state_S80 , state_T07 , state_T08 , state_C82 , state_C109 , state_P60 , state_B89 , state_P63 , state_B92 , state_L27 , state_S93 , state_B96 , state_B101 , state_S97 , state_S122 , state_C100 , state_S115 , state_P58 , state_B130 , state_L28 , state_S105 , state_T11 , state_T12 , state_L29 , state_S83 , state_S90 , state_L30 , state_P64 , state_P65 , state_L32 , state_L33 , state_S110 , state_C95 , state_C114 , state_T13 , state_T14 , state_T15 , state_S119 , state_T17 , state_C118 , state_T19 , state_T20 , state_T21 , state_T22 , state_L34 , state_S135 , state_L35 , state_X50 , state_X51 , state_P70 , state_P71 , state_L37 , state_L38 , state_P68 , state_P69 , state_S139 , state_L40 , state_C104 , state_L41 , state_T23 , state_T24 , state_L42 , state_S131 , state_B133 , state_B145 , state_B143 , state_S86 , state_S146 , state_P72 , state_P73 , state_S144 , state_S102 , state_C138 : hex_char;
	signal cmd_R1_ne1 , cmd_R2_ne7 , cmd_R3_ne14 , cmd_R3_ne52 , cmd_R4_ne47 , cmd_R4_ne48 , cmd_R5_ne84 , cmd_R5_ne82 , cmd_R5_ne32 , cmd_R6_ne84 , cmd_R6_ne85 , cmd_R6_ne100 , cmd_R6_ne101 , cmd_R6_ne44 , cmd_R7_ne89 , cmd_R7_ne30 , cmd_R8_ne90 , cmd_R8_ne91 , cmd_R8_ne30 , cmd_R9_ne105 , cmd_R9_ne98 , cmd_R9_ne96 , cmd_R10_ne4 , cmd_R10_ne106 , cmd_R11_ne26 , cmd_R11_ne65 , cmd_R12_ne44 , cmd_R12_ne101 , cmd_R13_ne65 , cmd_R13_ne102 , cmd_R14_ne70 , cmd_R14_ne104 , cmd_R14_ne21 , cmd_R15_ne78 , cmd_R15_ne93 , cmd_R16_ne93 , cmd_R16_ne96 , cmd_R17_ne95 , cmd_R18_ne97 , cmd_R18_ne94 , cmd_R19_ne98 , cmd_R19_ne105 , cmd_R20_ne101 , cmd_R20_ne100 , cmd_R21_ne103 , cmd_R21_ne64 , cmd_R22_ne106 , cmd_R22_ne99 , cmd_R23_ne7 , cmd_R23_ne9 , cmd_R24_ne9 , cmd_R24_ne95 , cmd_R25_ne95 , cmd_R25_ne59 , cmd_R26_ne95 , cmd_R26_ne9 , cmd_R27_ne23 , cmd_R27_ne26 , cmd_R28_ne24 , cmd_R28_ne64 , cmd_R28_ne103 , cmd_R28_ne67 , cmd_R29_ne67 , cmd_R29_ne70 , cmd_R30_ne67 , cmd_R30_ne103 , cmd_R31_ne99 , cmd_R31_ne97 , cmd_R32_ne99 , cmd_R32_ne106 , cmd_R32_ne4 , cmd_R33_ne96 , cmd_R33_ne93 , cmd_R33_ne78 , cmd_R34_ne96 , cmd_R34_ne98 , cmd_R35_ne21 , cmd_R36_ne21 , cmd_R36_ne79 , cmd_R36_ne78 , cmd_R37_ne21 , cmd_R37_ne94 , cmd_R37_ne97 , cmd_R37_ne99 , cmd_R38_ne1 , cmd_R38_ne9 , cmd_R39_ne9 , cmd_R39_ne1 , cmd_R40_ne9 , cmd_R40_ne7 , cmd_R41_ne17 , cmd_R41_ne59 , cmd_R41_ne95 , cmd_R42_ne59 , cmd_R42_ne11 , cmd_R42_ne52 , cmd_R43_ne59 , cmd_R43_ne17 , cmd_R44_ne52 , cmd_R44_ne11 , cmd_R44_ne59 , cmd_R44_ne95 , cmd_R45_ne52 , cmd_R45_ne14 , cmd_R46_ne23 , cmd_R46_ne64 , cmd_R46_ne103 , cmd_R46_ne67 , cmd_R47_ne64 , cmd_R47_ne23 , cmd_R48_ne64 , cmd_R48_ne24 , cmd_R49_ne24 , cmd_R49_ne26 , cmd_R50_ne26 , cmd_R50_ne23 , cmd_R51_ne26 , cmd_R51_ne24 , cmd_R52_ne83 , cmd_R52_ne30 , cmd_R53_ne29 , cmd_R53_ne30 , cmd_R54_ne30 , cmd_R54_ne29 , cmd_R54_ne110 , cmd_R55_ne30 , cmd_R55_ne83 , cmd_R56_ne32 , cmd_R56_ne110 , cmd_R57_ne29 , cmd_R58_ne110 , cmd_R58_ne32 , cmd_R59_ne110 , cmd_R59_ne29 , cmd_R60_ne102 , cmd_R60_ne44 , cmd_R61_ne44 , cmd_R61_ne43 , cmd_R61_ne48 , cmd_R62_ne44 , cmd_R62_ne102 , cmd_R62_ne65 , cmd_R62_ne26 , cmd_R63_ne17 , cmd_R63_ne78 , cmd_R64_ne78 , cmd_R64_ne17 , cmd_R65_ne78 , cmd_R65_ne79 , cmd_R65_ne77 , cmd_R66_ne78 , cmd_R66_ne79 , cmd_R66_ne21 , cmd_R67_ne83 , cmd_R67_ne32 , cmd_R68_ne32 , cmd_R68_ne83 , cmd_R69_ne32 , cmd_R69_ne82 , cmd_R69_ne41 , cmd_R70_ne32 , cmd_R70_ne82 , cmd_R70_ne84 , cmd_R71_ne88 , cmd_R71_ne86 , cmd_R72_ne86 , cmd_R72_ne88 , cmd_R73_ne86 , cmd_R73_ne87 , cmd_R73_ne91 , cmd_R73_ne30 , cmd_R74_ne30 , cmd_R74_ne89 , cmd_R75_ne30 , cmd_R75_ne91 , cmd_R75_ne87 , cmd_R75_ne86 , cmd_R76_ne30 , cmd_R76_ne91 , cmd_R76_ne90 , cmd_R77_ne41 , cmd_R77_ne82 , cmd_R77_ne32 , cmd_R78_ne41 , cmd_R78_ne85 , cmd_R78_ne100 , cmd_R78_ne101 , cmd_R78_ne44 , cmd_R79_ne85 , cmd_R79_ne41 , cmd_R80_ne85 , cmd_R80_ne84 , cmd_R81_ne77 , cmd_R81_ne52 , cmd_R82_ne94 , cmd_R82_ne77 , cmd_R83_ne94 , cmd_R83_ne21 , cmd_R84_ne110 , cmd_R84_ne100 , cmd_R84_ne101 , cmd_R84_ne44 , cmd_R85_ne100 , cmd_R85_ne110 , cmd_R86_ne100 , cmd_R86_ne85 , cmd_R87_ne104 , cmd_R87_ne70 , cmd_R88_ne21 , cmd_R88_ne104 , cmd_R89_ne77 , cmd_R89_ne79 , cmd_R89_ne78 , cmd_R90_ne77 , cmd_R90_ne94 , cmd_R90_ne97 , cmd_R90_ne99 , cmd_R91_ne52 , cmd_R91_ne77 : routeCommands := RELEASE;
	signal state_ne1 , state_ne4 , state_ne7 , state_ne9 , state_ne11 , state_ne14 , state_ne17 , state_ne23 , state_ne24 , state_ne26 , state_ne29 , state_ne30 , state_ne32 , state_ne41 , state_ne43 , state_ne44 , state_ne47 , state_ne48 , state_ne59 , state_ne64 , state_ne65 , state_ne67 , state_ne70 , state_ne78 , state_ne79 , state_ne82 , state_ne83 , state_ne84 , state_ne86 , state_ne87 , state_ne88 , state_ne89 , state_ne90 , state_ne91 , state_ne93 , state_ne94 , state_ne95 , state_ne96 , state_ne97 , state_ne98 , state_ne99 , state_ne100 , state_ne101 , state_ne102 , state_ne103 , state_ne105 , state_ne106 , state_ne85 , state_ne77 , state_ne104 , state_ne52 , state_ne21 , state_ne110 : hex_char;
	signal cmd_R25_Lc01 , cmd_R26_Lc01 , cmd_R41_Lc01 , cmd_R44_Lc01 : routeCommands := RELEASE;
	signal cmd_R23_68W02 , cmd_R38_68W02 , cmd_R39_68W02 , cmd_R40_68W02 , cmd_R1_68W02 , cmd_R2_68W02 , cmd_R26_68W02 , cmd_R41_69W03 , cmd_R42_69W03 , cmd_R43_69W03 , cmd_R44_69W03 , cmd_R64_69W03 , cmd_R25_69W03 , cmd_R81_69W03 , cmd_R3_69W04 , cmd_R42_69W04 , cmd_R44_69W04 , cmd_R45_69W04 , cmd_R25_69W04 , cmd_R81_69W04 , cmd_R36_Sw06 , cmd_R63_Sw06 , cmd_R64_Sw06 , cmd_R65_Sw06 , cmd_R66_Sw06 , cmd_R89_Sw06 , cmd_R43_Sw06 , cmd_R14_Sw06 , cmd_R33_Sw06 , cmd_R91_Sw06 , cmd_R47_70W01 , cmd_R48_70W01 , cmd_R21_70W01 , cmd_R27_70W02 , cmd_R49_70W02 , cmd_R50_70W02 , cmd_R51_70W02 , cmd_R62_70W02 , cmd_R47_70W02 , cmd_R48_70W02 , cmd_R52_Sw08 , cmd_R53_Sw08 , cmd_R54_Sw08 , cmd_R55_Sw08 , cmd_R57_Sw08 , cmd_R68_Sw08 , cmd_R73_Sw08 , cmd_R7_Sw08 , cmd_R8_Sw08 , cmd_R54_Sw09 , cmd_R56_Sw09 , cmd_R58_Sw09 , cmd_R59_Sw09 , cmd_R77_Sw09 , cmd_R67_Sw09 , cmd_R5_Sw09 , cmd_R73_Sw09 , cmd_R7_Sw09 , cmd_R8_Sw09 , cmd_R85_Sw09 , cmd_R7_Sw12 , cmd_R8_Sw12 , cmd_R73_Sw12 , cmd_R74_Sw12 , cmd_R75_Sw12 , cmd_R76_Sw12 , cmd_R53_Sw12 , cmd_R52_Sw12 , cmd_R5_Sw04 , cmd_R67_Sw04 , cmd_R68_Sw04 , cmd_R69_Sw04 , cmd_R70_Sw04 , cmd_R77_Sw04 , cmd_R55_Sw04 , cmd_R58_Sw04 , cmd_R60_71W01 , cmd_R61_71W01 , cmd_R62_71W01 , cmd_R78_71W01 , cmd_R13_71W01 , cmd_R6_71W01 , cmd_R84_71W01 , cmd_R4_71W02 , cmd_R61_71W02 , cmd_R78_71W02 , cmd_R6_71W02 , cmd_R84_71W02 , cmd_R71_Sw11 , cmd_R72_Sw11 , cmd_R73_Sw11 , cmd_R75_Sw11 , cmd_R8_Sw13 , cmd_R73_Sw13 , cmd_R75_Sw13 , cmd_R76_Sw13 , cmd_R6_Sw41 , cmd_R78_Sw41 , cmd_R84_Sw41 , cmd_R85_Sw41 , cmd_R86_Sw41 , cmd_R54_Sw41 , cmd_R56_Sw41 , cmd_R20_Sw41 : routeCommands := RELEASE;
	signal cmd_R5_Sw05 , cmd_R6_Sw05 , cmd_R69_Sw05 , cmd_R70_Sw05 , cmd_R77_Sw05 , cmd_R78_Sw05 , cmd_R79_Sw05 , cmd_R80_Sw05 , cmd_R36_Sw07 , cmd_R37_Sw07 , cmd_R65_Sw07 , cmd_R66_Sw07 , cmd_R82_Sw07 , cmd_R83_Sw07 , cmd_R89_Sw07 , cmd_R90_Sw07 : routeCommands := RELEASE;
	signal cmd_R14_Sw03 , cmd_R81_Sw03 , cmd_R88_Sw03 , cmd_R91_Sw03 : routeCommands := RELEASE;
	signal cmd_R1_T02 , cmd_R2_T06 , cmd_R3_T08 , cmd_R4_T12 , cmd_R5_T14 , cmd_R6_T14 , cmd_R7_T20 , cmd_R8_T22 , cmd_R9_T24 , cmd_R10_L25 , cmd_R11_L27 , cmd_R12_L28 , cmd_R13_L30 , cmd_R14_L32 , cmd_R15_L33 , cmd_R16_L34 , cmd_R17_L35 , cmd_R18_L37 , cmd_R19_L38 , cmd_R20_L40 , cmd_R21_L41 , cmd_R22_L42 , cmd_R23_J43 , cmd_R24_J46 , cmd_R25_X50 , cmd_R26_X51 , cmd_R27_P60 , cmd_R28_P63 , cmd_R29_P64 , cmd_R30_P65 , cmd_R31_P68 , cmd_R32_P69 , cmd_R33_P70 , cmd_R34_P71 , cmd_R35_P72 , cmd_R36_P73 , cmd_R37_P73 , cmd_R38_C78 , cmd_R39_S80 , cmd_R40_S80 , cmd_R41_C82 , cmd_R42_S83 , cmd_R43_S83 , cmd_R44_S86 , cmd_R45_S86 , cmd_R46_B89 , cmd_R47_S90 , cmd_R48_S90 , cmd_R49_B92 , cmd_R50_S93 , cmd_R51_S93 , cmd_R52_C95 , cmd_R53_B96 , cmd_R54_S97 , cmd_R55_S97 , cmd_R56_C100 , cmd_R57_B101 , cmd_R58_S102 , cmd_R59_S102 , cmd_R60_C104 , cmd_R61_S105 , cmd_R62_S105 , cmd_R63_C109 , cmd_R64_S110 , cmd_R65_S110 , cmd_R66_S110 , cmd_R67_C114 , cmd_R68_S115 , cmd_R69_S115 , cmd_R70_S115 , cmd_R71_C118 , cmd_R72_S119 , cmd_R73_S119 , cmd_R74_S122 , cmd_R75_S122 , cmd_R76_S122 , cmd_R77_B130 , cmd_R78_B130 , cmd_R79_S131 , cmd_R80_S131 , cmd_R81_B133 , cmd_R82_S135 , cmd_R83_S135 , cmd_R84_C138 , cmd_R85_S139 , cmd_R86_S139 , cmd_R87_B143 , cmd_R88_S144 , cmd_R89_B145 , cmd_R90_B145 , cmd_R91_S146 : routeCommands := RELEASE;
	signal cmd_R1_C78 , cmd_R2_J43 , cmd_R3_S146 , cmd_R4_L29 , cmd_R5_C100 , cmd_R6_S105 , cmd_R7_S97 , cmd_R8_S97 , cmd_R9_P70 , cmd_R10_L42 , cmd_R11_L30 , cmd_R12_L40 , cmd_R13_C104 , cmd_R14_P73 , cmd_R15_L34 , cmd_R16_P71 , cmd_R17_X50 , cmd_R18_S135 , cmd_R19_T23 , cmd_R20_S139 , cmd_R21_S90 , cmd_R22_P68 , cmd_R23_J46 , cmd_R24_L35 , cmd_R25_S83 , cmd_R26_S80 , cmd_R27_L27 , cmd_R28_P64 , cmd_R29_L32 , cmd_R30_L41 , cmd_R31_L37 , cmd_R32_T03 , cmd_R33_S110 , cmd_R34_L38 , cmd_R35_S144 , cmd_R36_L33 , cmd_R37_P69 , cmd_R38_J46 , cmd_R39_T01 , cmd_R40_T05 , cmd_R41_X51 , cmd_R42_S146 , cmd_R43_C109 , cmd_R44_X51 , cmd_R45_T07 , cmd_R46_P64 , cmd_R47_P60 , cmd_R48_B92 , cmd_R49_L27 , cmd_R50_B89 , cmd_R51_P63 , cmd_R52_S122 , cmd_R53_S122 , cmd_R54_C138 , cmd_R55_C114 , cmd_R56_C138 , cmd_R57_B96 , cmd_R58_S115 , cmd_R59_B101 , cmd_R60_L28 , cmd_R61_L29 , cmd_R62_S93 , cmd_R63_L33 , cmd_R64_C82 , cmd_R65_B133 , cmd_R66_P72 , cmd_R67_C100 , cmd_R68_C95 , cmd_R69_P58 , cmd_R70_T13 , cmd_R71_T15 , cmd_R72_T17 , cmd_R73_S97 , cmd_R74_T19 , cmd_R75_T15 , cmd_R76_T21 , cmd_R77_C100 , cmd_R78_S105 , cmd_R79_P58 , cmd_R80_T13 , cmd_R81_S86 , cmd_R82_B133 , cmd_R83_P72 , cmd_R84_S105 , cmd_R85_S102 , cmd_R86_S131 , cmd_R87_L32 , cmd_R88_B143 , cmd_R89_L33 , cmd_R90_P69 , cmd_R91_B145 : routeCommands := RELEASE;
begin
	levelCrossing_Lc01 : levelCrossing_0 port map(track_ne95 => tracks_i(36), track_ne9 => tracks_i(3), track_ne59 => tracks_i(18), R25_command => cmd_R25_Lc01, R26_command => cmd_R26_Lc01, R41_command => cmd_R41_Lc01, R44_command => cmd_R44_Lc01, indication => levelCrossings_i, command  => levelCrossings_o, correspondence => state_Lc01, clock => clock, reset => reset);
	singleSwitch_68W02 : singleSwitch_0 port map(R23_command => cmd_R23_68W02, R38_command => cmd_R38_68W02, R39_command => cmd_R39_68W02, R40_command => cmd_R40_68W02, R1_command => cmd_R1_68W02, R2_command => cmd_R2_68W02, R26_command => cmd_R26_68W02, indication => singleSwitches_i(0), command => singleSwitches_o(0), correspondence => state_68W02, clock => clock, reset => reset);
	singleSwitch_69W03 : singleSwitch_1 port map(R41_command => cmd_R41_69W03, R42_command => cmd_R42_69W03, R43_command => cmd_R43_69W03, R44_command => cmd_R44_69W03, R64_command => cmd_R64_69W03, R25_command => cmd_R25_69W03, R81_command => cmd_R81_69W03, indication => singleSwitches_i(1), command => singleSwitches_o(1), correspondence => state_69W03, clock => clock, reset => reset);
	singleSwitch_69W04 : singleSwitch_2 port map(R3_command => cmd_R3_69W04, R42_command => cmd_R42_69W04, R44_command => cmd_R44_69W04, R45_command => cmd_R45_69W04, R25_command => cmd_R25_69W04, R81_command => cmd_R81_69W04, indication => singleSwitches_i(2), command => singleSwitches_o(2), correspondence => state_69W04, clock => clock, reset => reset);
	singleSwitch_Sw06 : singleSwitch_3 port map(R36_command => cmd_R36_Sw06, R63_command => cmd_R63_Sw06, R64_command => cmd_R64_Sw06, R65_command => cmd_R65_Sw06, R66_command => cmd_R66_Sw06, R89_command => cmd_R89_Sw06, R43_command => cmd_R43_Sw06, R14_command => cmd_R14_Sw06, R33_command => cmd_R33_Sw06, R91_command => cmd_R91_Sw06, indication => singleSwitches_i(3), command => singleSwitches_o(3), correspondence => state_Sw06, clock => clock, reset => reset);
	singleSwitch_70W01 : singleSwitch_4 port map(R47_command => cmd_R47_70W01, R48_command => cmd_R48_70W01, R21_command => cmd_R21_70W01, indication => singleSwitches_i(4), command => singleSwitches_o(4), correspondence => state_70W01, clock => clock, reset => reset);
	singleSwitch_70W02 : singleSwitch_5 port map(R27_command => cmd_R27_70W02, R49_command => cmd_R49_70W02, R50_command => cmd_R50_70W02, R51_command => cmd_R51_70W02, R62_command => cmd_R62_70W02, R47_command => cmd_R47_70W02, R48_command => cmd_R48_70W02, indication => singleSwitches_i(5), command => singleSwitches_o(5), correspondence => state_70W02, clock => clock, reset => reset);
	singleSwitch_Sw08 : singleSwitch_6 port map(R52_command => cmd_R52_Sw08, R53_command => cmd_R53_Sw08, R54_command => cmd_R54_Sw08, R55_command => cmd_R55_Sw08, R57_command => cmd_R57_Sw08, R68_command => cmd_R68_Sw08, R73_command => cmd_R73_Sw08, R7_command => cmd_R7_Sw08, R8_command => cmd_R8_Sw08, indication => singleSwitches_i(6), command => singleSwitches_o(6), correspondence => state_Sw08, clock => clock, reset => reset);
	singleSwitch_Sw09 : singleSwitch_7 port map(R54_command => cmd_R54_Sw09, R56_command => cmd_R56_Sw09, R58_command => cmd_R58_Sw09, R59_command => cmd_R59_Sw09, R77_command => cmd_R77_Sw09, R67_command => cmd_R67_Sw09, R5_command => cmd_R5_Sw09, R73_command => cmd_R73_Sw09, R7_command => cmd_R7_Sw09, R8_command => cmd_R8_Sw09, R85_command => cmd_R85_Sw09, indication => singleSwitches_i(7), command => singleSwitches_o(7), correspondence => state_Sw09, clock => clock, reset => reset);
	singleSwitch_Sw12 : singleSwitch_8 port map(R7_command => cmd_R7_Sw12, R8_command => cmd_R8_Sw12, R73_command => cmd_R73_Sw12, R74_command => cmd_R74_Sw12, R75_command => cmd_R75_Sw12, R76_command => cmd_R76_Sw12, R53_command => cmd_R53_Sw12, R52_command => cmd_R52_Sw12, indication => singleSwitches_i(8), command => singleSwitches_o(8), correspondence => state_Sw12, clock => clock, reset => reset);
	singleSwitch_Sw04 : singleSwitch_9 port map(R5_command => cmd_R5_Sw04, R67_command => cmd_R67_Sw04, R68_command => cmd_R68_Sw04, R69_command => cmd_R69_Sw04, R70_command => cmd_R70_Sw04, R77_command => cmd_R77_Sw04, R55_command => cmd_R55_Sw04, R58_command => cmd_R58_Sw04, indication => singleSwitches_i(9), command => singleSwitches_o(9), correspondence => state_Sw04, clock => clock, reset => reset);
	singleSwitch_71W01 : singleSwitch_10 port map(R60_command => cmd_R60_71W01, R61_command => cmd_R61_71W01, R62_command => cmd_R62_71W01, R78_command => cmd_R78_71W01, R13_command => cmd_R13_71W01, R6_command => cmd_R6_71W01, R84_command => cmd_R84_71W01, indication => singleSwitches_i(10), command => singleSwitches_o(10), correspondence => state_71W01, clock => clock, reset => reset);
	singleSwitch_71W02 : singleSwitch_11 port map(R4_command => cmd_R4_71W02, R61_command => cmd_R61_71W02, R78_command => cmd_R78_71W02, R6_command => cmd_R6_71W02, R84_command => cmd_R84_71W02, indication => singleSwitches_i(11), command => singleSwitches_o(11), correspondence => state_71W02, clock => clock, reset => reset);
	singleSwitch_Sw11 : singleSwitch_12 port map(R71_command => cmd_R71_Sw11, R72_command => cmd_R72_Sw11, R73_command => cmd_R73_Sw11, R75_command => cmd_R75_Sw11, indication => singleSwitches_i(12), command => singleSwitches_o(12), correspondence => state_Sw11, clock => clock, reset => reset);
	singleSwitch_Sw13 : singleSwitch_13 port map(R8_command => cmd_R8_Sw13, R73_command => cmd_R73_Sw13, R75_command => cmd_R75_Sw13, R76_command => cmd_R76_Sw13, indication => singleSwitches_i(13), command => singleSwitches_o(13), correspondence => state_Sw13, clock => clock, reset => reset);
	singleSwitch_Sw41 : singleSwitch_14 port map(R6_command => cmd_R6_Sw41, R78_command => cmd_R78_Sw41, R84_command => cmd_R84_Sw41, R85_command => cmd_R85_Sw41, R86_command => cmd_R86_Sw41, R54_command => cmd_R54_Sw41, R56_command => cmd_R56_Sw41, R20_command => cmd_R20_Sw41, indication => singleSwitches_i(14), command => singleSwitches_o(14), correspondence => state_Sw41, clock => clock, reset => reset);
	scissorCrossing_Sw03 : scissorCrossing_0 port map(R14_command => cmd_R14_Sw03, R81_command => cmd_R81_Sw03, R88_command => cmd_R88_Sw03, R91_command => cmd_R91_Sw03, indication => scissorCrossings_i, command => scissorCrossings_o, correspondence => state_Sw03, clock => clock, reset => reset);
	doubleSwitch_Sw05 : doubleSwitch_0 port map(R5_command => cmd_R5_Sw05, R6_command => cmd_R6_Sw05, R69_command => cmd_R69_Sw05, R70_command => cmd_R70_Sw05, R77_command => cmd_R77_Sw05, R78_command => cmd_R78_Sw05, R79_command => cmd_R79_Sw05, R80_command => cmd_R80_Sw05, indication => doubleSwitches_i(0), command => doubleSwitches_o(0),correspondence=> state_Sw05, clock => clock, reset => reset);
	doubleSwitch_Sw07 : doubleSwitch_1 port map(R36_command => cmd_R36_Sw07, R37_command => cmd_R37_Sw07, R65_command => cmd_R65_Sw07, R66_command => cmd_R66_Sw07, R82_command => cmd_R82_Sw07, R83_command => cmd_R83_Sw07, R89_command => cmd_R89_Sw07, R90_command => cmd_R90_Sw07, indication => doubleSwitches_i(1), command => doubleSwitches_o(1),correspondence=> state_Sw07, clock => clock, reset => reset);
	railwaySignal_T01 : railwaySignal_0 port map(R39_command => cmd_R39_T01, track_ne1 => tracks_i(0), indication => signals_i(0), command => signals_o(0), correspondence_T01 => state_T01, clock => clock, reset => reset);
	railwaySignal_T02 : railwaySignal_1 port map(R1_command => cmd_R1_T02, track_ne1 => tracks_i(0), track_ne9 => tracks_i(3), correspondence_C78 => state_C78, correspondence_J46 => state_J46, s68W02_state => state_68W02, indication => signals_i(1), command => signals_o(1), correspondence_T02 => state_T02, clock => clock, reset => reset);
	railwaySignal_C78 : railwaySignal_2 port map(R38_command => cmd_R38_C78, R1_command => cmd_R1_C78, track_ne1 => tracks_i(0), track_ne9 => tracks_i(3), track_ne95 => tracks_i(36), correspondence_J46 => state_J46, correspondence_L35 => state_L35, s68W02_state => state_68W02, indication => signals_i(2), command => signals_o(2), correspondence_C78 => state_C78, clock => clock, reset => reset);
	railwaySignal_T03 : railwaySignal_3 port map(R32_command => cmd_R32_T03, track_ne4 => tracks_i(1), indication => signals_i(3), command => signals_o(3), correspondence_T03 => state_T03, clock => clock, reset => reset);
	railwaySignal_L25 : railwaySignal_4 port map(R10_command => cmd_R10_L25, track_ne4 => tracks_i(1), track_ne106 => tracks_i(46), track_ne99 => tracks_i(40), correspondence_L42 => state_L42, correspondence_P68 => state_P68, indication => signals_i(4), command => signals_o(4), correspondence_L25 => state_L25, clock => clock, reset => reset);
	railwaySignal_T05 : railwaySignal_5 port map(R40_command => cmd_R40_T05, track_ne7 => tracks_i(2), indication => signals_i(5), command => signals_o(5), correspondence_T05 => state_T05, clock => clock, reset => reset);
	railwaySignal_T06 : railwaySignal_6 port map(R2_command => cmd_R2_T06, track_ne7 => tracks_i(2), track_ne9 => tracks_i(3), correspondence_J43 => state_J43, correspondence_J46 => state_J46, s68W02_state => state_68W02, indication => signals_i(6), command => signals_o(6), correspondence_T06 => state_T06, clock => clock, reset => reset);
	railwaySignal_J43 : railwaySignal_7 port map(R23_command => cmd_R23_J43, R2_command => cmd_R2_J43, track_ne7 => tracks_i(2), track_ne9 => tracks_i(3), track_ne95 => tracks_i(36), correspondence_J46 => state_J46, correspondence_L35 => state_L35, s68W02_state => state_68W02, indication => signals_i(7), command => signals_o(7), correspondence_J43 => state_J43, clock => clock, reset => reset);
	railwaySignal_J46 : railwaySignal_8 port map(R24_command => cmd_R24_J46, R23_command => cmd_R23_J46, R38_command => cmd_R38_J46, track_ne9 => tracks_i(3), track_ne95 => tracks_i(36), correspondence_L35 => state_L35, correspondence_X50 => state_X50, indication => signals_i(8), command => signals_o(8), correspondence_J46 => state_J46, clock => clock, reset => reset);
	railwaySignal_S80 : railwaySignal_9 port map(R39_command => cmd_R39_S80, R40_command => cmd_R40_S80, R26_command => cmd_R26_S80, track_ne9 => tracks_i(3), track_ne1 => tracks_i(0), track_ne7 => tracks_i(2), correspondence_T01 => state_T01, correspondence_T05 => state_T05, s68W02_state => state_68W02, indication => signals_i(9), command => signals_o(9), correspondence_S80 => state_S80, clock => clock, reset => reset);
	railwaySignal_T07 : railwaySignal_10 port map(R45_command => cmd_R45_T07, track_ne14 => tracks_i(5), indication => signals_i(10), command => signals_o(10), correspondence_T07 => state_T07, clock => clock, reset => reset);
	railwaySignal_T08 : railwaySignal_11 port map(R3_command => cmd_R3_T08, track_ne14 => tracks_i(5), track_ne52 => tracks_i(50), track_ne77 => tracks_i(48), correspondence_S146 => state_S146, correspondence_B145 => state_B145, s69W04_state => state_69W04, Sw03_state => state_Sw03, indication => signals_i(11), command => signals_o(11), correspondence_T08 => state_T08, clock => clock, reset => reset);
	railwaySignal_C82 : railwaySignal_12 port map(R41_command => cmd_R41_C82, R64_command => cmd_R64_C82, track_ne17 => tracks_i(6), track_ne59 => tracks_i(18), track_ne95 => tracks_i(36), track_ne9 => tracks_i(3), correspondence_X51 => state_X51, correspondence_S80 => state_S80, s69W03_state => state_69W03, Lc01_state => state_Lc01, indication => signals_i(12), command => signals_o(12), correspondence_C82 => state_C82, clock => clock, reset => reset);
	railwaySignal_C109 : railwaySignal_13 port map(R63_command => cmd_R63_C109, R43_command => cmd_R43_C109, track_ne17 => tracks_i(6), track_ne78 => tracks_i(23), track_ne93 => tracks_i(34), correspondence_L33 => state_L33, correspondence_L34 => state_L34, Sw06_state => state_Sw06, indication => signals_i(13), command => signals_o(13), correspondence_C109 => state_C109, clock => clock, reset => reset);
	railwaySignal_P60 : railwaySignal_14 port map(R27_command => cmd_R27_P60, R47_command => cmd_R47_P60, track_ne23 => tracks_i(7), track_ne26 => tracks_i(9), track_ne65 => tracks_i(20), correspondence_L27 => state_L27, correspondence_L30 => state_L30, s70W02_state => state_70W02, indication => signals_i(14), command => signals_o(14), correspondence_P60 => state_P60, clock => clock, reset => reset);
	railwaySignal_B89 : railwaySignal_15 port map(R46_command => cmd_R46_B89, R50_command => cmd_R50_B89, track_ne23 => tracks_i(7), track_ne64 => tracks_i(19), track_ne103 => tracks_i(44), track_ne67 => tracks_i(21), track_ne70 => tracks_i(22), correspondence_P64 => state_P64, correspondence_L32 => state_L32, indication => signals_i(15), command => signals_o(15), correspondence_B89 => state_B89, clock => clock, reset => reset);
	railwaySignal_P63 : railwaySignal_16 port map(R28_command => cmd_R28_P63, R51_command => cmd_R51_P63, track_ne24 => tracks_i(8), track_ne64 => tracks_i(19), track_ne103 => tracks_i(44), track_ne67 => tracks_i(21), track_ne70 => tracks_i(22), correspondence_P64 => state_P64, correspondence_L32 => state_L32, indication => signals_i(16), command => signals_o(16), correspondence_P63 => state_P63, clock => clock, reset => reset);
	railwaySignal_B92 : railwaySignal_17 port map(R49_command => cmd_R49_B92, R48_command => cmd_R48_B92, track_ne24 => tracks_i(8), track_ne26 => tracks_i(9), track_ne65 => tracks_i(20), correspondence_L27 => state_L27, correspondence_L30 => state_L30, s70W02_state => state_70W02, indication => signals_i(17), command => signals_o(17), correspondence_B92 => state_B92, clock => clock, reset => reset);
	railwaySignal_L27 : railwaySignal_18 port map(R11_command => cmd_R11_L27, R27_command => cmd_R27_L27, R49_command => cmd_R49_L27, track_ne26 => tracks_i(9), track_ne65 => tracks_i(20), track_ne102 => tracks_i(43), correspondence_L30 => state_L30, correspondence_C104 => state_C104, indication => signals_i(18), command => signals_o(18), correspondence_L27 => state_L27, clock => clock, reset => reset);
	railwaySignal_S93 : railwaySignal_19 port map(R50_command => cmd_R50_S93, R51_command => cmd_R51_S93, R62_command => cmd_R62_S93, track_ne26 => tracks_i(9), track_ne23 => tracks_i(7), track_ne24 => tracks_i(8), track_ne67 => tracks_i(21), track_ne64 => tracks_i(19), track_ne103 => tracks_i(44), correspondence_B89 => state_B89, correspondence_P63 => state_P63, correspondence_P64 => state_P64, s70W02_state => state_70W02, indication => signals_i(19), command => signals_o(19), correspondence_S93 => state_S93, clock => clock, reset => reset);
	railwaySignal_B96 : railwaySignal_20 port map(R53_command => cmd_R53_B96, R57_command => cmd_R57_B96, track_ne29 => tracks_i(10), track_ne30 => tracks_i(11), track_ne87 => tracks_i(29), track_ne86 => tracks_i(28), track_ne91 => tracks_i(33), track_ne89 => tracks_i(31), track_ne90 => tracks_i(32), correspondence_S122 => state_S122, correspondence_T19 => state_T19, correspondence_T15 => state_T15, correspondence_T21 => state_T21, Sw08_state => state_Sw08, Sw12_state => state_Sw12, Sw11_state => state_Sw11, Sw13_state => state_Sw13, indication => signals_i(20), command => signals_o(20), correspondence_B96 => state_B96, clock => clock, reset => reset);
	railwaySignal_B101 : railwaySignal_21 port map(R57_command => cmd_R57_B101, R59_command => cmd_R59_B101, track_ne29 => tracks_i(10), track_ne30 => tracks_i(11), correspondence_B96 => state_B96, correspondence_S122 => state_S122, Sw08_state => state_Sw08, indication => signals_i(21), command => signals_o(21), correspondence_B101 => state_B101, clock => clock, reset => reset);
	railwaySignal_S97 : railwaySignal_22 port map(R54_command => cmd_R54_S97, R55_command => cmd_R55_S97, R7_command => cmd_R7_S97, R8_command => cmd_R8_S97, R73_command => cmd_R73_S97, track_ne30 => tracks_i(11), track_ne29 => tracks_i(10), track_ne110 => tracks_i(52), track_ne83 => tracks_i(26), track_ne100 => tracks_i(41), track_ne101 => tracks_i(42), track_ne44 => tracks_i(15), track_ne32 => tracks_i(12), correspondence_C138 => state_C138, correspondence_C114 => state_C114, correspondence_S105 => state_S105, correspondence_C100 => state_C100, Sw08_state => state_Sw08, Sw09_state => state_Sw09, Sw41_state => state_Sw41, Sw04_state => state_Sw04, indication => signals_i(22), command => signals_o(22), correspondence_S97 => state_S97, clock => clock, reset => reset);
	railwaySignal_S122 : railwaySignal_23 port map(R74_command => cmd_R74_S122, R75_command => cmd_R75_S122, R76_command => cmd_R76_S122, R52_command => cmd_R52_S122, R53_command => cmd_R53_S122, track_ne30 => tracks_i(11), track_ne89 => tracks_i(31), track_ne91 => tracks_i(33), track_ne87 => tracks_i(29), track_ne86 => tracks_i(28), track_ne90 => tracks_i(32), correspondence_T19 => state_T19, correspondence_T15 => state_T15, correspondence_T21 => state_T21, Sw12_state => state_Sw12, Sw11_state => state_Sw11, Sw13_state => state_Sw13, indication => signals_i(23), command => signals_o(23), correspondence_S122 => state_S122, clock => clock, reset => reset);
	railwaySignal_C100 : railwaySignal_24 port map(R56_command => cmd_R56_C100, R5_command => cmd_R5_C100, R67_command => cmd_R67_C100, R77_command => cmd_R77_C100, track_ne32 => tracks_i(12), track_ne110 => tracks_i(52), track_ne100 => tracks_i(41), track_ne101 => tracks_i(42), track_ne44 => tracks_i(15), correspondence_C138 => state_C138, correspondence_S105 => state_S105, Sw09_state => state_Sw09, Sw41_state => state_Sw41, indication => signals_i(24), command => signals_o(24), correspondence_C100 => state_C100, clock => clock, reset => reset);
	railwaySignal_S115 : railwaySignal_25 port map(R68_command => cmd_R68_S115, R69_command => cmd_R69_S115, R70_command => cmd_R70_S115, R58_command => cmd_R58_S115, track_ne32 => tracks_i(12), track_ne83 => tracks_i(26), track_ne82 => tracks_i(25), track_ne41 => tracks_i(13), track_ne84 => tracks_i(27), track_ne30 => tracks_i(11), correspondence_C95 => state_C95, correspondence_P58 => state_P58, correspondence_T13 => state_T13, correspondence_S122 => state_S122, Sw04_state => state_Sw04, Sw08_state => state_Sw08, Sw05_state => state_Sw05, indication => signals_i(25), command => signals_o(25), correspondence_S115 => state_S115, clock => clock, reset => reset);
	railwaySignal_P58 : railwaySignal_26 port map(R69_command => cmd_R69_P58, R79_command => cmd_R79_P58, track_ne41 => tracks_i(13), indication => signals_i(26), command => signals_o(26), correspondence_P58 => state_P58, clock => clock, reset => reset);
	railwaySignal_B130 : railwaySignal_27 port map(R77_command => cmd_R77_B130, R78_command => cmd_R78_B130, track_ne41 => tracks_i(13), track_ne82 => tracks_i(25), track_ne32 => tracks_i(12), track_ne85 => tracks_i(47), track_ne100 => tracks_i(41), track_ne101 => tracks_i(42), track_ne44 => tracks_i(15), track_ne110 => tracks_i(52), track_ne26 => tracks_i(9), track_ne43 => tracks_i(14), track_ne102 => tracks_i(43), track_ne48 => tracks_i(17), track_ne65 => tracks_i(20), correspondence_C100 => state_C100, correspondence_S105 => state_S105, correspondence_C138 => state_C138, correspondence_L29 => state_L29, correspondence_S93 => state_S93, Sw04_state => state_Sw04, Sw05_state => state_Sw05, Sw09_state => state_Sw09, Sw41_state => state_Sw41, s71W01_state => state_71W01, s71W02_state => state_71W02, indication => signals_i(27), command => signals_o(27), correspondence_B130 => state_B130, clock => clock, reset => reset);
	railwaySignal_L28 : railwaySignal_28 port map(R12_command => cmd_R12_L28, R60_command => cmd_R60_L28, track_ne44 => tracks_i(15), track_ne101 => tracks_i(42), track_ne100 => tracks_i(41), correspondence_L40 => state_L40, correspondence_S139 => state_S139, indication => signals_i(28), command => signals_o(28), correspondence_L28 => state_L28, clock => clock, reset => reset);
	railwaySignal_S105 : railwaySignal_29 port map(R61_command => cmd_R61_S105, R62_command => cmd_R62_S105, R6_command => cmd_R6_S105, R78_command => cmd_R78_S105, R84_command => cmd_R84_S105, track_ne44 => tracks_i(15), track_ne43 => tracks_i(14), track_ne48 => tracks_i(17), track_ne102 => tracks_i(43), track_ne65 => tracks_i(20), track_ne26 => tracks_i(9), track_ne23 => tracks_i(7), track_ne24 => tracks_i(8), correspondence_L29 => state_L29, correspondence_S93 => state_S93, correspondence_B89 => state_B89, correspondence_P63 => state_P63, s71W01_state => state_71W01, s71W02_state => state_71W02, s70W02_state => state_70W02, indication => signals_i(29), command => signals_o(29), correspondence_S105 => state_S105, clock => clock, reset => reset);
	railwaySignal_T11 : railwaySignal_30 port map(track_ne47 => tracks_i(16), indication => signals_i(30), command => signals_o(30), correspondence_T11 => state_T11, clock => clock, reset => reset);
	railwaySignal_T12 : railwaySignal_31 port map(R4_command => cmd_R4_T12, track_ne47 => tracks_i(16), track_ne48 => tracks_i(17), correspondence_L29 => state_L29, s71W02_state => state_71W02, indication => signals_i(31), command => signals_o(31), correspondence_T12 => state_T12, clock => clock, reset => reset);
	railwaySignal_L29 : railwaySignal_32 port map(R4_command => cmd_R4_L29, R61_command => cmd_R61_L29, track_ne48 => tracks_i(17), indication => signals_i(32), command => signals_o(32), correspondence_L29 => state_L29, clock => clock, reset => reset);
	railwaySignal_S83 : railwaySignal_33 port map(R42_command => cmd_R42_S83, R43_command => cmd_R43_S83, R25_command => cmd_R25_S83, track_ne59 => tracks_i(18), track_ne11 => tracks_i(4), track_ne52 => tracks_i(50), track_ne17 => tracks_i(6), track_ne77 => tracks_i(48), track_ne78 => tracks_i(23), correspondence_S146 => state_S146, correspondence_C109 => state_C109, correspondence_B145 => state_B145, correspondence_L33 => state_L33, s69W03_state => state_69W03, s69W04_state => state_69W04, Sw03_state => state_Sw03, Sw06_state => state_Sw06, indication => signals_i(33), command => signals_o(33), correspondence_S83 => state_S83, clock => clock, reset => reset);
	railwaySignal_S90 : railwaySignal_34 port map(R47_command => cmd_R47_S90, R48_command => cmd_R48_S90, R21_command => cmd_R21_S90, track_ne64 => tracks_i(19), track_ne23 => tracks_i(7), track_ne24 => tracks_i(8), track_ne26 => tracks_i(9), correspondence_P60 => state_P60, correspondence_B92 => state_B92, correspondence_L27 => state_L27, s70W01_state => state_70W01, s70W02_state => state_70W02, indication => signals_i(34), command => signals_o(34), correspondence_S90 => state_S90, clock => clock, reset => reset);
	railwaySignal_L30 : railwaySignal_35 port map(R13_command => cmd_R13_L30, R11_command => cmd_R11_L30, track_ne65 => tracks_i(20), track_ne102 => tracks_i(43), track_ne44 => tracks_i(15), correspondence_C104 => state_C104, correspondence_L28 => state_L28, s71W01_state => state_71W01, indication => signals_i(35), command => signals_o(35), correspondence_L30 => state_L30, clock => clock, reset => reset);
	railwaySignal_P64 : railwaySignal_36 port map(R29_command => cmd_R29_P64, R28_command => cmd_R28_P64, R46_command => cmd_R46_P64, track_ne67 => tracks_i(21), track_ne70 => tracks_i(22), track_ne104 => tracks_i(49), track_ne21 => tracks_i(51), correspondence_L32 => state_L32, correspondence_P73 => state_P73, Sw03_state => state_Sw03, indication => signals_i(36), command => signals_o(36), correspondence_P64 => state_P64, clock => clock, reset => reset);
	railwaySignal_P65 : railwaySignal_37 port map(R30_command => cmd_R30_P65, track_ne67 => tracks_i(21), track_ne103 => tracks_i(44), track_ne64 => tracks_i(19), correspondence_L41 => state_L41, correspondence_S90 => state_S90, indication => signals_i(37), command => signals_o(37), correspondence_P65 => state_P65, clock => clock, reset => reset);
	railwaySignal_L32 : railwaySignal_38 port map(R14_command => cmd_R14_L32, R29_command => cmd_R29_L32, R87_command => cmd_R87_L32, track_ne70 => tracks_i(22), track_ne104 => tracks_i(49), track_ne21 => tracks_i(51), track_ne97 => tracks_i(38), track_ne94 => tracks_i(35), track_ne79 => tracks_i(24), track_ne78 => tracks_i(23), track_ne99 => tracks_i(40), correspondence_P73 => state_P73, correspondence_L33 => state_L33, correspondence_P69 => state_P69, Sw03_state => state_Sw03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication => signals_i(38), command => signals_o(38), correspondence_L32 => state_L32, clock => clock, reset => reset);
	railwaySignal_L33 : railwaySignal_39 port map(R15_command => cmd_R15_L33, R36_command => cmd_R36_L33, R63_command => cmd_R63_L33, R89_command => cmd_R89_L33, track_ne78 => tracks_i(23), track_ne93 => tracks_i(34), track_ne96 => tracks_i(37), correspondence_L34 => state_L34, correspondence_P71 => state_P71, indication => signals_i(39), command => signals_o(39), correspondence_L33 => state_L33, clock => clock, reset => reset);
	railwaySignal_S110 : railwaySignal_40 port map(R64_command => cmd_R64_S110, R65_command => cmd_R65_S110, R66_command => cmd_R66_S110, R33_command => cmd_R33_S110, track_ne78 => tracks_i(23), track_ne17 => tracks_i(6), track_ne79 => tracks_i(24), track_ne77 => tracks_i(48), track_ne21 => tracks_i(51), track_ne59 => tracks_i(18), track_ne95 => tracks_i(36), track_ne52 => tracks_i(50), correspondence_C82 => state_C82, correspondence_B133 => state_B133, correspondence_P72 => state_P72, correspondence_X51 => state_X51, correspondence_S86 => state_S86, correspondence_S144 => state_S144, Sw06_state => state_Sw06, s69W03_state => state_69W03, Sw07_state => state_Sw07, Sw03_state => state_Sw03, indication => signals_i(40), command => signals_o(40), correspondence_S110 => state_S110, clock => clock, reset => reset);
	railwaySignal_C95 : railwaySignal_41 port map(R52_command => cmd_R52_C95, R68_command => cmd_R68_C95, track_ne83 => tracks_i(26), track_ne30 => tracks_i(11), track_ne87 => tracks_i(29), track_ne86 => tracks_i(28), track_ne91 => tracks_i(33), track_ne89 => tracks_i(31), track_ne90 => tracks_i(32), correspondence_S122 => state_S122, correspondence_T19 => state_T19, correspondence_T15 => state_T15, correspondence_T21 => state_T21, Sw08_state => state_Sw08, Sw12_state => state_Sw12, Sw11_state => state_Sw11, Sw13_state => state_Sw13, indication => signals_i(41), command => signals_o(41), correspondence_C95 => state_C95, clock => clock, reset => reset);
	railwaySignal_C114 : railwaySignal_42 port map(R67_command => cmd_R67_C114, R55_command => cmd_R55_C114, track_ne83 => tracks_i(26), track_ne32 => tracks_i(12), track_ne110 => tracks_i(52), correspondence_C100 => state_C100, correspondence_C138 => state_C138, Sw04_state => state_Sw04, Sw09_state => state_Sw09, indication => signals_i(42), command => signals_o(42), correspondence_C114 => state_C114, clock => clock, reset => reset);
	railwaySignal_T13 : railwaySignal_43 port map(R70_command => cmd_R70_T13, R80_command => cmd_R80_T13, track_ne84 => tracks_i(27), indication => signals_i(43), command => signals_o(43), correspondence_T13 => state_T13, clock => clock, reset => reset);
	railwaySignal_T14 : railwaySignal_44 port map(R5_command => cmd_R5_T14, R6_command => cmd_R6_T14, track_ne84 => tracks_i(27), track_ne82 => tracks_i(25), track_ne32 => tracks_i(12), track_ne85 => tracks_i(47), track_ne100 => tracks_i(41), track_ne101 => tracks_i(42), track_ne44 => tracks_i(15), track_ne110 => tracks_i(52), track_ne26 => tracks_i(9), track_ne43 => tracks_i(14), track_ne102 => tracks_i(43), track_ne48 => tracks_i(17), track_ne65 => tracks_i(20), correspondence_C100 => state_C100, correspondence_S105 => state_S105, correspondence_C138 => state_C138, correspondence_L29 => state_L29, correspondence_S93 => state_S93, Sw04_state => state_Sw04, Sw05_state => state_Sw05, Sw09_state => state_Sw09, Sw41_state => state_Sw41, s71W01_state => state_71W01, s71W02_state => state_71W02, indication => signals_i(44), command => signals_o(44), correspondence_T14 => state_T14, clock => clock, reset => reset);
	railwaySignal_T15 : railwaySignal_45 port map(R71_command => cmd_R71_T15, R75_command => cmd_R75_T15, track_ne86 => tracks_i(28), indication => signals_i(45), command => signals_o(45), correspondence_T15 => state_T15, clock => clock, reset => reset);
	railwaySignal_S119 : railwaySignal_46 port map(R72_command => cmd_R72_S119, R73_command => cmd_R73_S119, track_ne86 => tracks_i(28), track_ne88 => tracks_i(30), track_ne87 => tracks_i(29), track_ne91 => tracks_i(33), track_ne30 => tracks_i(11), track_ne83 => tracks_i(26), track_ne29 => tracks_i(10), track_ne110 => tracks_i(52), correspondence_T17 => state_T17, correspondence_S97 => state_S97, correspondence_C138 => state_C138, correspondence_C114 => state_C114, Sw11_state => state_Sw11, Sw12_state => state_Sw12, Sw13_state => state_Sw13, Sw08_state => state_Sw08, Sw09_state => state_Sw09, indication => signals_i(46), command => signals_o(46), correspondence_S119 => state_S119, clock => clock, reset => reset);
	railwaySignal_T17 : railwaySignal_47 port map(R72_command => cmd_R72_T17, track_ne88 => tracks_i(30), indication => signals_i(47), command => signals_o(47), correspondence_T17 => state_T17, clock => clock, reset => reset);
	railwaySignal_C118 : railwaySignal_48 port map(R71_command => cmd_R71_C118, track_ne88 => tracks_i(30), track_ne86 => tracks_i(28), correspondence_T15 => state_T15, Sw11_state => state_Sw11, indication => signals_i(48), command => signals_o(48), correspondence_C118 => state_C118, clock => clock, reset => reset);
	railwaySignal_T19 : railwaySignal_49 port map(R74_command => cmd_R74_T19, track_ne89 => tracks_i(31), indication => signals_i(49), command => signals_o(49), correspondence_T19 => state_T19, clock => clock, reset => reset);
	railwaySignal_T20 : railwaySignal_50 port map(R7_command => cmd_R7_T20, track_ne89 => tracks_i(31), track_ne30 => tracks_i(11), track_ne83 => tracks_i(26), track_ne29 => tracks_i(10), track_ne110 => tracks_i(52), correspondence_S97 => state_S97, correspondence_C138 => state_C138, correspondence_C114 => state_C114, Sw12_state => state_Sw12, Sw08_state => state_Sw08, Sw09_state => state_Sw09, indication => signals_i(50), command => signals_o(50), correspondence_T20 => state_T20, clock => clock, reset => reset);
	railwaySignal_T21 : railwaySignal_51 port map(R76_command => cmd_R76_T21, track_ne90 => tracks_i(32), indication => signals_i(51), command => signals_o(51), correspondence_T21 => state_T21, clock => clock, reset => reset);
	railwaySignal_T22 : railwaySignal_52 port map(R8_command => cmd_R8_T22, track_ne90 => tracks_i(32), track_ne91 => tracks_i(33), track_ne30 => tracks_i(11), track_ne83 => tracks_i(26), track_ne29 => tracks_i(10), track_ne110 => tracks_i(52), correspondence_S97 => state_S97, correspondence_C138 => state_C138, correspondence_C114 => state_C114, Sw12_state => state_Sw12, Sw13_state => state_Sw13, Sw08_state => state_Sw08, Sw09_state => state_Sw09, indication => signals_i(52), command => signals_o(52), correspondence_T22 => state_T22, clock => clock, reset => reset);
	railwaySignal_L34 : railwaySignal_53 port map(R16_command => cmd_R16_L34, R15_command => cmd_R15_L34, track_ne93 => tracks_i(34), track_ne96 => tracks_i(37), track_ne98 => tracks_i(39), correspondence_P71 => state_P71, correspondence_L38 => state_L38, indication => signals_i(53), command => signals_o(53), correspondence_L34 => state_L34, clock => clock, reset => reset);
	railwaySignal_S135 : railwaySignal_54 port map(R82_command => cmd_R82_S135, R83_command => cmd_R83_S135, R18_command => cmd_R18_S135, track_ne94 => tracks_i(35), track_ne77 => tracks_i(48), track_ne21 => tracks_i(51), track_ne52 => tracks_i(50), correspondence_B133 => state_B133, correspondence_P72 => state_P72, correspondence_S86 => state_S86, correspondence_S144 => state_S144, Sw07_state => state_Sw07, Sw03_state => state_Sw03, indication => signals_i(54), command => signals_o(54), correspondence_S135 => state_S135, clock => clock, reset => reset);
	railwaySignal_L35 : railwaySignal_55 port map(R17_command => cmd_R17_L35, R24_command => cmd_R24_L35, track_ne95 => tracks_i(36), track_ne59 => tracks_i(18), correspondence_X50 => state_X50, correspondence_S83 => state_S83, indication => signals_i(55), command => signals_o(55), correspondence_L35 => state_L35, clock => clock, reset => reset);
	railwaySignal_X50 : railwaySignal_56 port map(R25_command => cmd_R25_X50, R17_command => cmd_R17_X50, track_ne95 => tracks_i(36), track_ne59 => tracks_i(18), track_ne17 => tracks_i(6), track_ne11 => tracks_i(4), track_ne52 => tracks_i(50), correspondence_S83 => state_S83, correspondence_S146 => state_S146, correspondence_C109 => state_C109, s69W03_state => state_69W03, s69W04_state => state_69W04, Lc01_state => state_Lc01, indication => signals_i(56), command => signals_o(56), correspondence_X50 => state_X50, clock => clock, reset => reset);
	railwaySignal_X51 : railwaySignal_57 port map(R26_command => cmd_R26_X51, R41_command => cmd_R41_X51, R44_command => cmd_R44_X51, track_ne95 => tracks_i(36), track_ne9 => tracks_i(3), track_ne7 => tracks_i(2), track_ne1 => tracks_i(0), correspondence_S80 => state_S80, correspondence_T01 => state_T01, correspondence_T05 => state_T05, s68W02_state => state_68W02, Lc01_state => state_Lc01, indication => signals_i(57), command => signals_o(57), correspondence_X51 => state_X51, clock => clock, reset => reset);
	railwaySignal_P70 : railwaySignal_58 port map(R33_command => cmd_R33_P70, R9_command => cmd_R9_P70, track_ne96 => tracks_i(37), track_ne93 => tracks_i(34), track_ne78 => tracks_i(23), track_ne17 => tracks_i(6), track_ne79 => tracks_i(24), track_ne21 => tracks_i(51), track_ne77 => tracks_i(48), correspondence_S110 => state_S110, correspondence_C82 => state_C82, correspondence_B133 => state_B133, correspondence_P72 => state_P72, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication => signals_i(58), command => signals_o(58), correspondence_P70 => state_P70, clock => clock, reset => reset);
	railwaySignal_P71 : railwaySignal_59 port map(R34_command => cmd_R34_P71, R16_command => cmd_R16_P71, track_ne96 => tracks_i(37), track_ne98 => tracks_i(39), track_ne105 => tracks_i(45), correspondence_L38 => state_L38, correspondence_T23 => state_T23, indication => signals_i(59), command => signals_o(59), correspondence_P71 => state_P71, clock => clock, reset => reset);
	railwaySignal_L37 : railwaySignal_60 port map(R18_command => cmd_R18_L37, R31_command => cmd_R31_L37, track_ne97 => tracks_i(38), track_ne94 => tracks_i(35), track_ne21 => tracks_i(51), track_ne77 => tracks_i(48), correspondence_S135 => state_S135, correspondence_B133 => state_B133, correspondence_P72 => state_P72, Sw07_state => state_Sw07, indication => signals_i(60), command => signals_o(60), correspondence_L37 => state_L37, clock => clock, reset => reset);
	railwaySignal_L38 : railwaySignal_61 port map(R19_command => cmd_R19_L38, R34_command => cmd_R34_L38, track_ne98 => tracks_i(39), track_ne105 => tracks_i(45), correspondence_T23 => state_T23, indication => signals_i(61), command => signals_o(61), correspondence_L38 => state_L38, clock => clock, reset => reset);
	railwaySignal_P68 : railwaySignal_62 port map(R31_command => cmd_R31_P68, R22_command => cmd_R22_P68, track_ne99 => tracks_i(40), track_ne97 => tracks_i(38), track_ne94 => tracks_i(35), correspondence_L37 => state_L37, correspondence_S135 => state_S135, indication => signals_i(62), command => signals_o(62), correspondence_P68 => state_P68, clock => clock, reset => reset);
	railwaySignal_P69 : railwaySignal_63 port map(R32_command => cmd_R32_P69, R37_command => cmd_R37_P69, R90_command => cmd_R90_P69, track_ne99 => tracks_i(40), track_ne106 => tracks_i(46), track_ne4 => tracks_i(1), correspondence_T03 => state_T03, indication => signals_i(63), command => signals_o(63), correspondence_P69 => state_P69, clock => clock, reset => reset);
	railwaySignal_S139 : railwaySignal_64 port map(R85_command => cmd_R85_S139, R86_command => cmd_R86_S139, R20_command => cmd_R20_S139, track_ne100 => tracks_i(41), track_ne110 => tracks_i(52), track_ne85 => tracks_i(47), track_ne32 => tracks_i(12), track_ne29 => tracks_i(10), track_ne84 => tracks_i(27), track_ne41 => tracks_i(13), correspondence_S102 => state_S102, correspondence_S131 => state_S131, correspondence_S115 => state_S115, correspondence_B101 => state_B101, correspondence_P58 => state_P58, correspondence_T13 => state_T13, Sw41_state => state_Sw41, Sw09_state => state_Sw09, Sw05_state => state_Sw05, indication => signals_i(64), command => signals_o(64), correspondence_S139 => state_S139, clock => clock, reset => reset);
	railwaySignal_L40 : railwaySignal_65 port map(R20_command => cmd_R20_L40, R12_command => cmd_R12_L40, track_ne101 => tracks_i(42), track_ne100 => tracks_i(41), track_ne85 => tracks_i(47), track_ne110 => tracks_i(52), correspondence_S139 => state_S139, correspondence_S102 => state_S102, correspondence_S131 => state_S131, Sw41_state => state_Sw41, indication => signals_i(65), command => signals_o(65), correspondence_L40 => state_L40, clock => clock, reset => reset);
	railwaySignal_C104 : railwaySignal_66 port map(R60_command => cmd_R60_C104, R13_command => cmd_R13_C104, track_ne102 => tracks_i(43), track_ne44 => tracks_i(15), track_ne101 => tracks_i(42), correspondence_L28 => state_L28, correspondence_L40 => state_L40, s71W01_state => state_71W01, indication => signals_i(66), command => signals_o(66), correspondence_C104 => state_C104, clock => clock, reset => reset);
	railwaySignal_L41 : railwaySignal_67 port map(R21_command => cmd_R21_L41, R30_command => cmd_R30_L41, track_ne103 => tracks_i(44), track_ne64 => tracks_i(19), track_ne23 => tracks_i(7), track_ne24 => tracks_i(8), correspondence_S90 => state_S90, correspondence_P60 => state_P60, correspondence_B92 => state_B92, s70W01_state => state_70W01, indication => signals_i(67), command => signals_o(67), correspondence_L41 => state_L41, clock => clock, reset => reset);
	railwaySignal_T23 : railwaySignal_68 port map(R19_command => cmd_R19_T23, track_ne105 => tracks_i(45), indication => signals_i(68), command => signals_o(68), correspondence_T23 => state_T23, clock => clock, reset => reset);
	railwaySignal_T24 : railwaySignal_69 port map(R9_command => cmd_R9_T24, track_ne105 => tracks_i(45), track_ne98 => tracks_i(39), track_ne96 => tracks_i(37), track_ne93 => tracks_i(34), track_ne78 => tracks_i(23), correspondence_P70 => state_P70, correspondence_S110 => state_S110, indication => signals_i(69), command => signals_o(69), correspondence_T24 => state_T24, clock => clock, reset => reset);
	railwaySignal_L42 : railwaySignal_70 port map(R22_command => cmd_R22_L42, R10_command => cmd_R10_L42, track_ne106 => tracks_i(46), track_ne99 => tracks_i(40), track_ne97 => tracks_i(38), correspondence_P68 => state_P68, correspondence_L37 => state_L37, indication => signals_i(70), command => signals_o(70), correspondence_L42 => state_L42, clock => clock, reset => reset);
	railwaySignal_S131 : railwaySignal_71 port map(R79_command => cmd_R79_S131, R80_command => cmd_R80_S131, R86_command => cmd_R86_S131, track_ne85 => tracks_i(47), track_ne41 => tracks_i(13), track_ne84 => tracks_i(27), correspondence_P58 => state_P58, correspondence_T13 => state_T13, Sw05_state => state_Sw05, indication => signals_i(71), command => signals_o(71), correspondence_S131 => state_S131, clock => clock, reset => reset);
	railwaySignal_B133 : railwaySignal_72 port map(R81_command => cmd_R81_B133, R65_command => cmd_R65_B133, R82_command => cmd_R82_B133, track_ne77 => tracks_i(48), track_ne52 => tracks_i(50), track_ne59 => tracks_i(18), track_ne11 => tracks_i(4), track_ne14 => tracks_i(5), track_ne95 => tracks_i(36), correspondence_S86 => state_S86, correspondence_X51 => state_X51, correspondence_T07 => state_T07, Sw03_state => state_Sw03, s69W03_state => state_69W03, s69W04_state => state_69W04, indication => signals_i(72), command => signals_o(72), correspondence_B133 => state_B133, clock => clock, reset => reset);
	railwaySignal_B145 : railwaySignal_73 port map(R89_command => cmd_R89_B145, R90_command => cmd_R90_B145, R91_command => cmd_R91_B145, track_ne77 => tracks_i(48), track_ne79 => tracks_i(24), track_ne78 => tracks_i(23), track_ne94 => tracks_i(35), track_ne97 => tracks_i(38), track_ne99 => tracks_i(40), track_ne93 => tracks_i(34), track_ne4 => tracks_i(1), track_ne106 => tracks_i(46), correspondence_L33 => state_L33, correspondence_P69 => state_P69, correspondence_L34 => state_L34, correspondence_T03 => state_T03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication => signals_i(73), command => signals_o(73), correspondence_B145 => state_B145, clock => clock, reset => reset);
	railwaySignal_B143 : railwaySignal_74 port map(R87_command => cmd_R87_B143, R88_command => cmd_R88_B143, track_ne104 => tracks_i(49), track_ne70 => tracks_i(22), track_ne21 => tracks_i(51), correspondence_L32 => state_L32, correspondence_P73 => state_P73, Sw03_state => state_Sw03, indication => signals_i(74), command => signals_o(74), correspondence_B143 => state_B143, clock => clock, reset => reset);
	railwaySignal_S86 : railwaySignal_75 port map(R44_command => cmd_R44_S86, R45_command => cmd_R45_S86, R81_command => cmd_R81_S86, track_ne52 => tracks_i(50), track_ne11 => tracks_i(4), track_ne59 => tracks_i(18), track_ne95 => tracks_i(36), track_ne14 => tracks_i(5), track_ne9 => tracks_i(3), correspondence_X51 => state_X51, correspondence_T07 => state_T07, correspondence_S80 => state_S80, s69W03_state => state_69W03, s69W04_state => state_69W04, Lc01_state => state_Lc01, indication => signals_i(75), command => signals_o(75), correspondence_S86 => state_S86, clock => clock, reset => reset);
	railwaySignal_S146 : railwaySignal_76 port map(R91_command => cmd_R91_S146, R3_command => cmd_R3_S146, R42_command => cmd_R42_S146, track_ne52 => tracks_i(50), track_ne77 => tracks_i(48), track_ne97 => tracks_i(38), track_ne94 => tracks_i(35), track_ne79 => tracks_i(24), track_ne78 => tracks_i(23), track_ne99 => tracks_i(40), correspondence_B145 => state_B145, correspondence_L33 => state_L33, correspondence_P69 => state_P69, Sw03_state => state_Sw03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication => signals_i(76), command => signals_o(76), correspondence_S146 => state_S146, clock => clock, reset => reset);
	railwaySignal_P72 : railwaySignal_77 port map(R35_command => cmd_R35_P72, R66_command => cmd_R66_P72, R83_command => cmd_R83_P72, track_ne21 => tracks_i(51), track_ne104 => tracks_i(49), correspondence_S144 => state_S144, correspondence_B143 => state_B143, Sw03_state => state_Sw03, indication => signals_i(77), command => signals_o(77), correspondence_P72 => state_P72, clock => clock, reset => reset);
	railwaySignal_P73 : railwaySignal_78 port map(R36_command => cmd_R36_P73, R37_command => cmd_R37_P73, R14_command => cmd_R14_P73, track_ne21 => tracks_i(51), track_ne79 => tracks_i(24), track_ne78 => tracks_i(23), track_ne94 => tracks_i(35), track_ne97 => tracks_i(38), track_ne99 => tracks_i(40), track_ne93 => tracks_i(34), track_ne4 => tracks_i(1), track_ne106 => tracks_i(46), correspondence_L33 => state_L33, correspondence_P69 => state_P69, correspondence_L34 => state_L34, correspondence_T03 => state_T03, Sw06_state => state_Sw06, Sw07_state => state_Sw07, indication => signals_i(78), command => signals_o(78), correspondence_P73 => state_P73, clock => clock, reset => reset);
	railwaySignal_S144 : railwaySignal_79 port map(R88_command => cmd_R88_S144, R35_command => cmd_R35_S144, track_ne21 => tracks_i(51), track_ne104 => tracks_i(49), track_ne70 => tracks_i(22), correspondence_B143 => state_B143, correspondence_L32 => state_L32, Sw03_state => state_Sw03, indication => signals_i(79), command => signals_o(79), correspondence_S144 => state_S144, clock => clock, reset => reset);
	railwaySignal_S102 : railwaySignal_80 port map(R58_command => cmd_R58_S102, R59_command => cmd_R59_S102, R85_command => cmd_R85_S102, track_ne110 => tracks_i(52), track_ne32 => tracks_i(12), track_ne29 => tracks_i(10), track_ne84 => tracks_i(27), track_ne83 => tracks_i(26), track_ne41 => tracks_i(13), track_ne82 => tracks_i(25), correspondence_S115 => state_S115, correspondence_B101 => state_B101, correspondence_C95 => state_C95, correspondence_P58 => state_P58, correspondence_T13 => state_T13, correspondence_B96 => state_B96, Sw09_state => state_Sw09, Sw04_state => state_Sw04, Sw05_state => state_Sw05, indication => signals_i(80), command => signals_o(80), correspondence_S102 => state_S102, clock => clock, reset => reset);
	railwaySignal_C138 : railwaySignal_81 port map(R84_command => cmd_R84_C138, R54_command => cmd_R54_C138, R56_command => cmd_R56_C138, track_ne110 => tracks_i(52), track_ne100 => tracks_i(41), track_ne101 => tracks_i(42), track_ne44 => tracks_i(15), track_ne26 => tracks_i(9), track_ne43 => tracks_i(14), track_ne102 => tracks_i(43), track_ne48 => tracks_i(17), track_ne65 => tracks_i(20), correspondence_S105 => state_S105, correspondence_L29 => state_L29, correspondence_S93 => state_S93, Sw41_state => state_Sw41, s71W01_state => state_71W01, s71W02_state => state_71W02, indication => signals_i(81), command => signals_o(81), correspondence_C138 => state_C138, clock => clock, reset => reset);
	node_ne1 : node_0 port map(track_i => tracks_i(0), track_o => state_ne1, R1_command => cmd_R1_ne1, R38_command => cmd_R38_ne1, R39_command => cmd_R39_ne1, reset => reset);
	node_ne4 : node_1 port map(track_i => tracks_i(1), track_o => state_ne4, R10_command => cmd_R10_ne4, R32_command => cmd_R32_ne4, reset => reset);
	node_ne7 : node_2 port map(track_i => tracks_i(2), track_o => state_ne7, R2_command => cmd_R2_ne7, R23_command => cmd_R23_ne7, R40_command => cmd_R40_ne7, reset => reset);
	node_ne9 : node_3 port map(track_i => tracks_i(3), track_o => state_ne9, R23_command => cmd_R23_ne9, R24_command => cmd_R24_ne9, R26_command => cmd_R26_ne9, R38_command => cmd_R38_ne9, R39_command => cmd_R39_ne9, R40_command => cmd_R40_ne9, reset => reset);
	node_ne11 : node_4 port map(track_i => tracks_i(4), track_o => state_ne11, R42_command => cmd_R42_ne11, R44_command => cmd_R44_ne11, reset => reset);
	node_ne14 : node_5 port map(track_i => tracks_i(5), track_o => state_ne14, R3_command => cmd_R3_ne14, R45_command => cmd_R45_ne14, reset => reset);
	node_ne17 : node_6 port map(track_i => tracks_i(6), track_o => state_ne17, R41_command => cmd_R41_ne17, R43_command => cmd_R43_ne17, R63_command => cmd_R63_ne17, R64_command => cmd_R64_ne17, reset => reset);
	node_ne23 : node_7 port map(track_i => tracks_i(7), track_o => state_ne23, R27_command => cmd_R27_ne23, R46_command => cmd_R46_ne23, R47_command => cmd_R47_ne23, R50_command => cmd_R50_ne23, reset => reset);
	node_ne24 : node_8 port map(track_i => tracks_i(8), track_o => state_ne24, R28_command => cmd_R28_ne24, R48_command => cmd_R48_ne24, R49_command => cmd_R49_ne24, R51_command => cmd_R51_ne24, reset => reset);
	node_ne26 : node_9 port map(track_i => tracks_i(9), track_o => state_ne26, R11_command => cmd_R11_ne26, R27_command => cmd_R27_ne26, R49_command => cmd_R49_ne26, R50_command => cmd_R50_ne26, R51_command => cmd_R51_ne26, R62_command => cmd_R62_ne26, reset => reset);
	node_ne29 : node_10 port map(track_i => tracks_i(10), track_o => state_ne29, R53_command => cmd_R53_ne29, R54_command => cmd_R54_ne29, R57_command => cmd_R57_ne29, R59_command => cmd_R59_ne29, reset => reset);
	node_ne30 : node_11 port map(track_i => tracks_i(11), track_o => state_ne30, R7_command => cmd_R7_ne30, R8_command => cmd_R8_ne30, R52_command => cmd_R52_ne30, R53_command => cmd_R53_ne30, R54_command => cmd_R54_ne30, R55_command => cmd_R55_ne30, R73_command => cmd_R73_ne30, R74_command => cmd_R74_ne30, R75_command => cmd_R75_ne30, R76_command => cmd_R76_ne30, reset => reset);
	node_ne32 : node_12 port map(track_i => tracks_i(12), track_o => state_ne32, R5_command => cmd_R5_ne32, R56_command => cmd_R56_ne32, R58_command => cmd_R58_ne32, R67_command => cmd_R67_ne32, R68_command => cmd_R68_ne32, R69_command => cmd_R69_ne32, R70_command => cmd_R70_ne32, R77_command => cmd_R77_ne32, reset => reset);
	node_ne41 : node_13 port map(track_i => tracks_i(13), track_o => state_ne41, R69_command => cmd_R69_ne41, R77_command => cmd_R77_ne41, R78_command => cmd_R78_ne41, R79_command => cmd_R79_ne41, reset => reset);
	node_ne43 : node_14 port map(track_i => tracks_i(14), track_o => state_ne43, R61_command => cmd_R61_ne43, reset => reset);
	node_ne44 : node_15 port map(track_i => tracks_i(15), track_o => state_ne44, R6_command => cmd_R6_ne44, R12_command => cmd_R12_ne44, R60_command => cmd_R60_ne44, R61_command => cmd_R61_ne44, R62_command => cmd_R62_ne44, R78_command => cmd_R78_ne44, R84_command => cmd_R84_ne44, reset => reset);
	node_ne47 : node_16 port map(track_i => tracks_i(16), track_o => state_ne47, R4_command => cmd_R4_ne47, reset => reset);
	node_ne48 : node_17 port map(track_i => tracks_i(17), track_o => state_ne48, R4_command => cmd_R4_ne48, R61_command => cmd_R61_ne48, reset => reset);
	node_ne59 : node_18 port map(track_i => tracks_i(18), track_o => state_ne59, R25_command => cmd_R25_ne59, R41_command => cmd_R41_ne59, R42_command => cmd_R42_ne59, R43_command => cmd_R43_ne59, R44_command => cmd_R44_ne59, reset => reset);
	node_ne64 : node_19 port map(track_i => tracks_i(19), track_o => state_ne64, R21_command => cmd_R21_ne64, R28_command => cmd_R28_ne64, R46_command => cmd_R46_ne64, R47_command => cmd_R47_ne64, R48_command => cmd_R48_ne64, reset => reset);
	node_ne65 : node_20 port map(track_i => tracks_i(20), track_o => state_ne65, R11_command => cmd_R11_ne65, R13_command => cmd_R13_ne65, R62_command => cmd_R62_ne65, reset => reset);
	node_ne67 : node_21 port map(track_i => tracks_i(21), track_o => state_ne67, R28_command => cmd_R28_ne67, R29_command => cmd_R29_ne67, R30_command => cmd_R30_ne67, R46_command => cmd_R46_ne67, reset => reset);
	node_ne70 : node_22 port map(track_i => tracks_i(22), track_o => state_ne70, R14_command => cmd_R14_ne70, R29_command => cmd_R29_ne70, R87_command => cmd_R87_ne70, reset => reset);
	node_ne78 : node_23 port map(track_i => tracks_i(23), track_o => state_ne78, R15_command => cmd_R15_ne78, R33_command => cmd_R33_ne78, R36_command => cmd_R36_ne78, R63_command => cmd_R63_ne78, R64_command => cmd_R64_ne78, R65_command => cmd_R65_ne78, R66_command => cmd_R66_ne78, R89_command => cmd_R89_ne78, reset => reset);
	node_ne79 : node_24 port map(track_i => tracks_i(24), track_o => state_ne79, R36_command => cmd_R36_ne79, R65_command => cmd_R65_ne79, R66_command => cmd_R66_ne79, R89_command => cmd_R89_ne79, reset => reset);
	node_ne82 : node_25 port map(track_i => tracks_i(25), track_o => state_ne82, R5_command => cmd_R5_ne82, R69_command => cmd_R69_ne82, R70_command => cmd_R70_ne82, R77_command => cmd_R77_ne82, reset => reset);
	node_ne83 : node_26 port map(track_i => tracks_i(26), track_o => state_ne83, R52_command => cmd_R52_ne83, R55_command => cmd_R55_ne83, R67_command => cmd_R67_ne83, R68_command => cmd_R68_ne83, reset => reset);
	node_ne84 : node_27 port map(track_i => tracks_i(27), track_o => state_ne84, R5_command => cmd_R5_ne84, R6_command => cmd_R6_ne84, R70_command => cmd_R70_ne84, R80_command => cmd_R80_ne84, reset => reset);
	node_ne86 : node_28 port map(track_i => tracks_i(28), track_o => state_ne86, R71_command => cmd_R71_ne86, R72_command => cmd_R72_ne86, R73_command => cmd_R73_ne86, R75_command => cmd_R75_ne86, reset => reset);
	node_ne87 : node_29 port map(track_i => tracks_i(29), track_o => state_ne87, R73_command => cmd_R73_ne87, R75_command => cmd_R75_ne87, reset => reset);
	node_ne88 : node_30 port map(track_i => tracks_i(30), track_o => state_ne88, R71_command => cmd_R71_ne88, R72_command => cmd_R72_ne88, reset => reset);
	node_ne89 : node_31 port map(track_i => tracks_i(31), track_o => state_ne89, R7_command => cmd_R7_ne89, R74_command => cmd_R74_ne89, reset => reset);
	node_ne90 : node_32 port map(track_i => tracks_i(32), track_o => state_ne90, R8_command => cmd_R8_ne90, R76_command => cmd_R76_ne90, reset => reset);
	node_ne91 : node_33 port map(track_i => tracks_i(33), track_o => state_ne91, R8_command => cmd_R8_ne91, R73_command => cmd_R73_ne91, R75_command => cmd_R75_ne91, R76_command => cmd_R76_ne91, reset => reset);
	node_ne93 : node_34 port map(track_i => tracks_i(34), track_o => state_ne93, R15_command => cmd_R15_ne93, R16_command => cmd_R16_ne93, R33_command => cmd_R33_ne93, reset => reset);
	node_ne94 : node_35 port map(track_i => tracks_i(35), track_o => state_ne94, R18_command => cmd_R18_ne94, R37_command => cmd_R37_ne94, R82_command => cmd_R82_ne94, R83_command => cmd_R83_ne94, R90_command => cmd_R90_ne94, reset => reset);
	node_ne95 : node_36 port map(track_i => tracks_i(36), track_o => state_ne95, R17_command => cmd_R17_ne95, R24_command => cmd_R24_ne95, R25_command => cmd_R25_ne95, R26_command => cmd_R26_ne95, R41_command => cmd_R41_ne95, R44_command => cmd_R44_ne95, reset => reset);
	node_ne96 : node_37 port map(track_i => tracks_i(37), track_o => state_ne96, R9_command => cmd_R9_ne96, R16_command => cmd_R16_ne96, R33_command => cmd_R33_ne96, R34_command => cmd_R34_ne96, reset => reset);
	node_ne97 : node_38 port map(track_i => tracks_i(38), track_o => state_ne97, R18_command => cmd_R18_ne97, R31_command => cmd_R31_ne97, R37_command => cmd_R37_ne97, R90_command => cmd_R90_ne97, reset => reset);
	node_ne98 : node_39 port map(track_i => tracks_i(39), track_o => state_ne98, R9_command => cmd_R9_ne98, R19_command => cmd_R19_ne98, R34_command => cmd_R34_ne98, reset => reset);
	node_ne99 : node_40 port map(track_i => tracks_i(40), track_o => state_ne99, R22_command => cmd_R22_ne99, R31_command => cmd_R31_ne99, R32_command => cmd_R32_ne99, R37_command => cmd_R37_ne99, R90_command => cmd_R90_ne99, reset => reset);
	node_ne100 : node_41 port map(track_i => tracks_i(41), track_o => state_ne100, R6_command => cmd_R6_ne100, R20_command => cmd_R20_ne100, R78_command => cmd_R78_ne100, R84_command => cmd_R84_ne100, R85_command => cmd_R85_ne100, R86_command => cmd_R86_ne100, reset => reset);
	node_ne101 : node_42 port map(track_i => tracks_i(42), track_o => state_ne101, R6_command => cmd_R6_ne101, R12_command => cmd_R12_ne101, R20_command => cmd_R20_ne101, R78_command => cmd_R78_ne101, R84_command => cmd_R84_ne101, reset => reset);
	node_ne102 : node_43 port map(track_i => tracks_i(43), track_o => state_ne102, R13_command => cmd_R13_ne102, R60_command => cmd_R60_ne102, R62_command => cmd_R62_ne102, reset => reset);
	node_ne103 : node_44 port map(track_i => tracks_i(44), track_o => state_ne103, R21_command => cmd_R21_ne103, R28_command => cmd_R28_ne103, R30_command => cmd_R30_ne103, R46_command => cmd_R46_ne103, reset => reset);
	node_ne105 : node_45 port map(track_i => tracks_i(45), track_o => state_ne105, R9_command => cmd_R9_ne105, R19_command => cmd_R19_ne105, reset => reset);
	node_ne106 : node_46 port map(track_i => tracks_i(46), track_o => state_ne106, R10_command => cmd_R10_ne106, R22_command => cmd_R22_ne106, R32_command => cmd_R32_ne106, reset => reset);
	node_ne85 : node_47 port map(track_i => tracks_i(47), track_o => state_ne85, R6_command => cmd_R6_ne85, R78_command => cmd_R78_ne85, R79_command => cmd_R79_ne85, R80_command => cmd_R80_ne85, R86_command => cmd_R86_ne85, reset => reset);
	node_ne77 : node_48 port map(track_i => tracks_i(48), track_o => state_ne77, R65_command => cmd_R65_ne77, R81_command => cmd_R81_ne77, R82_command => cmd_R82_ne77, R89_command => cmd_R89_ne77, R90_command => cmd_R90_ne77, R91_command => cmd_R91_ne77, reset => reset);
	node_ne104 : node_49 port map(track_i => tracks_i(49), track_o => state_ne104, R14_command => cmd_R14_ne104, R87_command => cmd_R87_ne104, R88_command => cmd_R88_ne104, reset => reset);
	node_ne52 : node_50 port map(track_i => tracks_i(50), track_o => state_ne52, R3_command => cmd_R3_ne52, R42_command => cmd_R42_ne52, R44_command => cmd_R44_ne52, R45_command => cmd_R45_ne52, R81_command => cmd_R81_ne52, R91_command => cmd_R91_ne52, reset => reset);
	node_ne21 : node_51 port map(track_i => tracks_i(51), track_o => state_ne21, R14_command => cmd_R14_ne21, R35_command => cmd_R35_ne21, R36_command => cmd_R36_ne21, R37_command => cmd_R37_ne21, R66_command => cmd_R66_ne21, R83_command => cmd_R83_ne21, R88_command => cmd_R88_ne21, reset => reset);
	node_ne110 : node_52 port map(track_i => tracks_i(52), track_o => state_ne110, R54_command => cmd_R54_ne110, R56_command => cmd_R56_ne110, R58_command => cmd_R58_ne110, R59_command => cmd_R59_ne110, R84_command => cmd_R84_ne110, R85_command => cmd_R85_ne110, reset => reset);
	route_R1 : route_0 port map(routeRequest => routes_i(0), ne1_command => cmd_R1_ne1, track_ne1 => state_ne1, s68W02_command => cmd_R1_68W02, s68W02_state => state_68W02, T02_state => state_T02, T02_command => cmd_R1_T02, C78_state => state_C78, C78_command =>cmd_R1_C78, routeExecute => routes_o(0), clock => clock, reset => reset);
	route_R2 : route_1 port map(routeRequest => routes_i(1), ne7_command => cmd_R2_ne7, track_ne7 => state_ne7, s68W02_command => cmd_R2_68W02, s68W02_state => state_68W02, T06_state => state_T06, T06_command => cmd_R2_T06, J43_state => state_J43, J43_command =>cmd_R2_J43, routeExecute => routes_o(1), clock => clock, reset => reset);
	route_R3 : route_2 port map(routeRequest => routes_i(2), ne14_command => cmd_R3_ne14, track_ne14 => state_ne14, ne52_command => cmd_R3_ne52, track_ne52 => state_ne52, s69W04_command => cmd_R3_69W04, s69W04_state => state_69W04, T08_state => state_T08, T08_command => cmd_R3_T08, S146_state => state_S146, S146_command =>cmd_R3_S146, routeExecute => routes_o(2), clock => clock, reset => reset);
	route_R4 : route_3 port map(routeRequest => routes_i(3), ne47_command => cmd_R4_ne47, track_ne47 => state_ne47, ne48_command => cmd_R4_ne48, track_ne48 => state_ne48, s71W02_command => cmd_R4_71W02, s71W02_state => state_71W02, T12_state => state_T12, T12_command => cmd_R4_T12, L29_state => state_L29, L29_command =>cmd_R4_L29, routeExecute => routes_o(3), clock => clock, reset => reset);
	route_R5 : route_4 port map(routeRequest => routes_i(4), ne32_command => cmd_R5_ne32, track_ne32 => state_ne32, ne82_command => cmd_R5_ne82, track_ne82 => state_ne82, ne84_command => cmd_R5_ne84, track_ne84 => state_ne84, Sw09_command => cmd_R5_Sw09, Sw09_state => state_Sw09, Sw04_command => cmd_R5_Sw04, Sw04_state => state_Sw04, Sw05_command => cmd_R5_Sw05, Sw05_state => state_Sw05, T14_state => state_T14, T14_command => cmd_R5_T14, C100_state => state_C100, C100_command =>cmd_R5_C100, routeExecute => routes_o(4), clock => clock, reset => reset);
	route_R6 : route_5 port map(routeRequest => routes_i(5), ne44_command => cmd_R6_ne44, track_ne44 => state_ne44, ne84_command => cmd_R6_ne84, track_ne84 => state_ne84, ne100_command => cmd_R6_ne100, track_ne100 => state_ne100, ne101_command => cmd_R6_ne101, track_ne101 => state_ne101, ne85_command => cmd_R6_ne85, track_ne85 => state_ne85, s71W01_command => cmd_R6_71W01, s71W01_state => state_71W01, s71W02_command => cmd_R6_71W02, s71W02_state => state_71W02, Sw41_command => cmd_R6_Sw41, Sw41_state => state_Sw41, Sw05_command => cmd_R6_Sw05, Sw05_state => state_Sw05, T14_state => state_T14, T14_command => cmd_R6_T14, S105_state => state_S105, S105_command =>cmd_R6_S105, routeExecute => routes_o(5), clock => clock, reset => reset);
	route_R7 : route_6 port map(routeRequest => routes_i(6), ne30_command => cmd_R7_ne30, track_ne30 => state_ne30, ne89_command => cmd_R7_ne89, track_ne89 => state_ne89, Sw08_command => cmd_R7_Sw08, Sw08_state => state_Sw08, Sw09_command => cmd_R7_Sw09, Sw09_state => state_Sw09, Sw12_command => cmd_R7_Sw12, Sw12_state => state_Sw12, T20_state => state_T20, T20_command => cmd_R7_T20, S97_state => state_S97, S97_command =>cmd_R7_S97, routeExecute => routes_o(6), clock => clock, reset => reset);
	route_R8 : route_7 port map(routeRequest => routes_i(7), ne30_command => cmd_R8_ne30, track_ne30 => state_ne30, ne90_command => cmd_R8_ne90, track_ne90 => state_ne90, ne91_command => cmd_R8_ne91, track_ne91 => state_ne91, Sw08_command => cmd_R8_Sw08, Sw08_state => state_Sw08, Sw09_command => cmd_R8_Sw09, Sw09_state => state_Sw09, Sw12_command => cmd_R8_Sw12, Sw12_state => state_Sw12, Sw13_command => cmd_R8_Sw13, Sw13_state => state_Sw13, T22_state => state_T22, T22_command => cmd_R8_T22, S97_state => state_S97, S97_command =>cmd_R8_S97, routeExecute => routes_o(7), clock => clock, reset => reset);
	route_R9 : route_8 port map(routeRequest => routes_i(8), ne96_command => cmd_R9_ne96, track_ne96 => state_ne96, ne98_command => cmd_R9_ne98, track_ne98 => state_ne98, ne105_command => cmd_R9_ne105, track_ne105 => state_ne105, T24_state => state_T24, T24_command => cmd_R9_T24, P70_state => state_P70, P70_command =>cmd_R9_P70, routeExecute => routes_o(8), clock => clock, reset => reset);
	route_R10 : route_9 port map(routeRequest => routes_i(9), ne4_command => cmd_R10_ne4, track_ne4 => state_ne4, ne106_command => cmd_R10_ne106, track_ne106 => state_ne106, L25_state => state_L25, L25_command => cmd_R10_L25, L42_state => state_L42, L42_command =>cmd_R10_L42, routeExecute => routes_o(9), clock => clock, reset => reset);
	route_R11 : route_10 port map(routeRequest => routes_i(10), ne26_command => cmd_R11_ne26, track_ne26 => state_ne26, ne65_command => cmd_R11_ne65, track_ne65 => state_ne65, L27_state => state_L27, L27_command => cmd_R11_L27, L30_state => state_L30, L30_command =>cmd_R11_L30, routeExecute => routes_o(10), clock => clock, reset => reset);
	route_R12 : route_11 port map(routeRequest => routes_i(11), ne44_command => cmd_R12_ne44, track_ne44 => state_ne44, ne101_command => cmd_R12_ne101, track_ne101 => state_ne101, L28_state => state_L28, L28_command => cmd_R12_L28, L40_state => state_L40, L40_command =>cmd_R12_L40, routeExecute => routes_o(11), clock => clock, reset => reset);
	route_R13 : route_12 port map(routeRequest => routes_i(12), ne65_command => cmd_R13_ne65, track_ne65 => state_ne65, ne102_command => cmd_R13_ne102, track_ne102 => state_ne102, s71W01_command => cmd_R13_71W01, s71W01_state => state_71W01, L30_state => state_L30, L30_command => cmd_R13_L30, C104_state => state_C104, C104_command =>cmd_R13_C104, routeExecute => routes_o(12), clock => clock, reset => reset);
	route_R14 : route_13 port map(routeRequest => routes_i(13), ne70_command => cmd_R14_ne70, track_ne70 => state_ne70, ne104_command => cmd_R14_ne104, track_ne104 => state_ne104, ne21_command => cmd_R14_ne21, track_ne21 => state_ne21, Sw06_command => cmd_R14_Sw06, Sw06_state => state_Sw06, Sw03_command => cmd_R14_Sw03, Sw03_state => state_Sw03, L32_state => state_L32, L32_command => cmd_R14_L32, P73_state => state_P73, P73_command =>cmd_R14_P73, routeExecute => routes_o(13), clock => clock, reset => reset);
	route_R15 : route_14 port map(routeRequest => routes_i(14), ne78_command => cmd_R15_ne78, track_ne78 => state_ne78, ne93_command => cmd_R15_ne93, track_ne93 => state_ne93, L33_state => state_L33, L33_command => cmd_R15_L33, L34_state => state_L34, L34_command =>cmd_R15_L34, routeExecute => routes_o(14), clock => clock, reset => reset);
	route_R16 : route_15 port map(routeRequest => routes_i(15), ne93_command => cmd_R16_ne93, track_ne93 => state_ne93, ne96_command => cmd_R16_ne96, track_ne96 => state_ne96, L34_state => state_L34, L34_command => cmd_R16_L34, P71_state => state_P71, P71_command =>cmd_R16_P71, routeExecute => routes_o(15), clock => clock, reset => reset);
	route_R17 : route_16 port map(routeRequest => routes_i(16), ne95_command => cmd_R17_ne95, track_ne95 => state_ne95, L35_state => state_L35, L35_command => cmd_R17_L35, X50_state => state_X50, X50_command =>cmd_R17_X50, routeExecute => routes_o(16), clock => clock, reset => reset);
	route_R18 : route_17 port map(routeRequest => routes_i(17), ne94_command => cmd_R18_ne94, track_ne94 => state_ne94, ne97_command => cmd_R18_ne97, track_ne97 => state_ne97, L37_state => state_L37, L37_command => cmd_R18_L37, S135_state => state_S135, S135_command =>cmd_R18_S135, routeExecute => routes_o(17), clock => clock, reset => reset);
	route_R19 : route_18 port map(routeRequest => routes_i(18), ne98_command => cmd_R19_ne98, track_ne98 => state_ne98, ne105_command => cmd_R19_ne105, track_ne105 => state_ne105, L38_state => state_L38, L38_command => cmd_R19_L38, T23_state => state_T23, T23_command =>cmd_R19_T23, routeExecute => routes_o(18), clock => clock, reset => reset);
	route_R20 : route_19 port map(routeRequest => routes_i(19), ne100_command => cmd_R20_ne100, track_ne100 => state_ne100, ne101_command => cmd_R20_ne101, track_ne101 => state_ne101, Sw41_command => cmd_R20_Sw41, Sw41_state => state_Sw41, L40_state => state_L40, L40_command => cmd_R20_L40, S139_state => state_S139, S139_command =>cmd_R20_S139, routeExecute => routes_o(19), clock => clock, reset => reset);
	route_R21 : route_20 port map(routeRequest => routes_i(20), ne64_command => cmd_R21_ne64, track_ne64 => state_ne64, ne103_command => cmd_R21_ne103, track_ne103 => state_ne103, s70W01_command => cmd_R21_70W01, s70W01_state => state_70W01, L41_state => state_L41, L41_command => cmd_R21_L41, S90_state => state_S90, S90_command =>cmd_R21_S90, routeExecute => routes_o(20), clock => clock, reset => reset);
	route_R22 : route_21 port map(routeRequest => routes_i(21), ne99_command => cmd_R22_ne99, track_ne99 => state_ne99, ne106_command => cmd_R22_ne106, track_ne106 => state_ne106, L42_state => state_L42, L42_command => cmd_R22_L42, P68_state => state_P68, P68_command =>cmd_R22_P68, routeExecute => routes_o(21), clock => clock, reset => reset);
	route_R23 : route_22 port map(routeRequest => routes_i(22), ne7_command => cmd_R23_ne7, track_ne7 => state_ne7, ne9_command => cmd_R23_ne9, track_ne9 => state_ne9, s68W02_command => cmd_R23_68W02, s68W02_state => state_68W02, J43_state => state_J43, J43_command => cmd_R23_J43, J46_state => state_J46, J46_command =>cmd_R23_J46, routeExecute => routes_o(22), clock => clock, reset => reset);
	route_R24 : route_23 port map(routeRequest => routes_i(23), ne9_command => cmd_R24_ne9, track_ne9 => state_ne9, ne95_command => cmd_R24_ne95, track_ne95 => state_ne95, J46_state => state_J46, J46_command => cmd_R24_J46, L35_state => state_L35, L35_command =>cmd_R24_L35, routeExecute => routes_o(23), clock => clock, reset => reset);
	route_R25 : route_24 port map(routeRequest => routes_i(24), ne59_command => cmd_R25_ne59, track_ne59 => state_ne59, ne95_command => cmd_R25_ne95, track_ne95 => state_ne95, Lc01_command => cmd_R25_Lc01, Lc01_state => state_Lc01, s69W03_command => cmd_R25_69W03, s69W03_state => state_69W03, s69W04_command => cmd_R25_69W04, s69W04_state => state_69W04, X50_state => state_X50, X50_command => cmd_R25_X50, S83_state => state_S83, S83_command =>cmd_R25_S83, routeExecute => routes_o(24), clock => clock, reset => reset);
	route_R26 : route_25 port map(routeRequest => routes_i(25), ne9_command => cmd_R26_ne9, track_ne9 => state_ne9, ne95_command => cmd_R26_ne95, track_ne95 => state_ne95, Lc01_command => cmd_R26_Lc01, Lc01_state => state_Lc01, s68W02_command => cmd_R26_68W02, s68W02_state => state_68W02, X51_state => state_X51, X51_command => cmd_R26_X51, S80_state => state_S80, S80_command =>cmd_R26_S80, routeExecute => routes_o(25), clock => clock, reset => reset);
	route_R27 : route_26 port map(routeRequest => routes_i(26), ne23_command => cmd_R27_ne23, track_ne23 => state_ne23, ne26_command => cmd_R27_ne26, track_ne26 => state_ne26, s70W02_command => cmd_R27_70W02, s70W02_state => state_70W02, P60_state => state_P60, P60_command => cmd_R27_P60, L27_state => state_L27, L27_command =>cmd_R27_L27, routeExecute => routes_o(26), clock => clock, reset => reset);
	route_R28 : route_27 port map(routeRequest => routes_i(27), ne24_command => cmd_R28_ne24, track_ne24 => state_ne24, ne64_command => cmd_R28_ne64, track_ne64 => state_ne64, ne67_command => cmd_R28_ne67, track_ne67 => state_ne67, ne103_command => cmd_R28_ne103, track_ne103 => state_ne103, P63_state => state_P63, P63_command => cmd_R28_P63, P64_state => state_P64, P64_command =>cmd_R28_P64, routeExecute => routes_o(27), clock => clock, reset => reset);
	route_R29 : route_28 port map(routeRequest => routes_i(28), ne67_command => cmd_R29_ne67, track_ne67 => state_ne67, ne70_command => cmd_R29_ne70, track_ne70 => state_ne70, P64_state => state_P64, P64_command => cmd_R29_P64, L32_state => state_L32, L32_command =>cmd_R29_L32, routeExecute => routes_o(28), clock => clock, reset => reset);
	route_R30 : route_29 port map(routeRequest => routes_i(29), ne67_command => cmd_R30_ne67, track_ne67 => state_ne67, ne103_command => cmd_R30_ne103, track_ne103 => state_ne103, P65_state => state_P65, P65_command => cmd_R30_P65, L41_state => state_L41, L41_command =>cmd_R30_L41, routeExecute => routes_o(29), clock => clock, reset => reset);
	route_R31 : route_30 port map(routeRequest => routes_i(30), ne97_command => cmd_R31_ne97, track_ne97 => state_ne97, ne99_command => cmd_R31_ne99, track_ne99 => state_ne99, P68_state => state_P68, P68_command => cmd_R31_P68, L37_state => state_L37, L37_command =>cmd_R31_L37, routeExecute => routes_o(30), clock => clock, reset => reset);
	route_R32 : route_31 port map(routeRequest => routes_i(31), ne4_command => cmd_R32_ne4, track_ne4 => state_ne4, ne99_command => cmd_R32_ne99, track_ne99 => state_ne99, ne106_command => cmd_R32_ne106, track_ne106 => state_ne106, P69_state => state_P69, P69_command => cmd_R32_P69, T03_state => state_T03, T03_command =>cmd_R32_T03, routeExecute => routes_o(31), clock => clock, reset => reset);
	route_R33 : route_32 port map(routeRequest => routes_i(32), ne78_command => cmd_R33_ne78, track_ne78 => state_ne78, ne93_command => cmd_R33_ne93, track_ne93 => state_ne93, ne96_command => cmd_R33_ne96, track_ne96 => state_ne96, Sw06_command => cmd_R33_Sw06, Sw06_state => state_Sw06, P70_state => state_P70, P70_command => cmd_R33_P70, S110_state => state_S110, S110_command =>cmd_R33_S110, routeExecute => routes_o(32), clock => clock, reset => reset);
	route_R34 : route_33 port map(routeRequest => routes_i(33), ne96_command => cmd_R34_ne96, track_ne96 => state_ne96, ne98_command => cmd_R34_ne98, track_ne98 => state_ne98, P71_state => state_P71, P71_command => cmd_R34_P71, L38_state => state_L38, L38_command =>cmd_R34_L38, routeExecute => routes_o(33), clock => clock, reset => reset);
	route_R35 : route_34 port map(routeRequest => routes_i(34), ne21_command => cmd_R35_ne21, track_ne21 => state_ne21, P72_state => state_P72, P72_command => cmd_R35_P72, S144_state => state_S144, S144_command =>cmd_R35_S144, routeExecute => routes_o(34), clock => clock, reset => reset);
	route_R36 : route_35 port map(routeRequest => routes_i(35), ne78_command => cmd_R36_ne78, track_ne78 => state_ne78, ne79_command => cmd_R36_ne79, track_ne79 => state_ne79, ne21_command => cmd_R36_ne21, track_ne21 => state_ne21, Sw06_command => cmd_R36_Sw06, Sw06_state => state_Sw06, Sw07_command => cmd_R36_Sw07, Sw07_state => state_Sw07, P73_state => state_P73, P73_command => cmd_R36_P73, L33_state => state_L33, L33_command =>cmd_R36_L33, routeExecute => routes_o(35), clock => clock, reset => reset);
	route_R37 : route_36 port map(routeRequest => routes_i(36), ne94_command => cmd_R37_ne94, track_ne94 => state_ne94, ne97_command => cmd_R37_ne97, track_ne97 => state_ne97, ne99_command => cmd_R37_ne99, track_ne99 => state_ne99, ne21_command => cmd_R37_ne21, track_ne21 => state_ne21, Sw07_command => cmd_R37_Sw07, Sw07_state => state_Sw07, P73_state => state_P73, P73_command => cmd_R37_P73, P69_state => state_P69, P69_command =>cmd_R37_P69, routeExecute => routes_o(36), clock => clock, reset => reset);
	route_R38 : route_37 port map(routeRequest => routes_i(37), ne1_command => cmd_R38_ne1, track_ne1 => state_ne1, ne9_command => cmd_R38_ne9, track_ne9 => state_ne9, s68W02_command => cmd_R38_68W02, s68W02_state => state_68W02, C78_state => state_C78, C78_command => cmd_R38_C78, J46_state => state_J46, J46_command =>cmd_R38_J46, routeExecute => routes_o(37), clock => clock, reset => reset);
	route_R39 : route_38 port map(routeRequest => routes_i(38), ne1_command => cmd_R39_ne1, track_ne1 => state_ne1, ne9_command => cmd_R39_ne9, track_ne9 => state_ne9, s68W02_command => cmd_R39_68W02, s68W02_state => state_68W02, S80_state => state_S80, S80_command => cmd_R39_S80, T01_state => state_T01, T01_command =>cmd_R39_T01, routeExecute => routes_o(38), clock => clock, reset => reset);
	route_R40 : route_39 port map(routeRequest => routes_i(39), ne7_command => cmd_R40_ne7, track_ne7 => state_ne7, ne9_command => cmd_R40_ne9, track_ne9 => state_ne9, s68W02_command => cmd_R40_68W02, s68W02_state => state_68W02, S80_state => state_S80, S80_command => cmd_R40_S80, T05_state => state_T05, T05_command =>cmd_R40_T05, routeExecute => routes_o(39), clock => clock, reset => reset);
	route_R41 : route_40 port map(routeRequest => routes_i(40), ne17_command => cmd_R41_ne17, track_ne17 => state_ne17, ne59_command => cmd_R41_ne59, track_ne59 => state_ne59, ne95_command => cmd_R41_ne95, track_ne95 => state_ne95, Lc01_command => cmd_R41_Lc01, Lc01_state => state_Lc01, s69W03_command => cmd_R41_69W03, s69W03_state => state_69W03, C82_state => state_C82, C82_command => cmd_R41_C82, X51_state => state_X51, X51_command =>cmd_R41_X51, routeExecute => routes_o(40), clock => clock, reset => reset);
	route_R42 : route_41 port map(routeRequest => routes_i(41), ne11_command => cmd_R42_ne11, track_ne11 => state_ne11, ne59_command => cmd_R42_ne59, track_ne59 => state_ne59, ne52_command => cmd_R42_ne52, track_ne52 => state_ne52, s69W03_command => cmd_R42_69W03, s69W03_state => state_69W03, s69W04_command => cmd_R42_69W04, s69W04_state => state_69W04, S83_state => state_S83, S83_command => cmd_R42_S83, S146_state => state_S146, S146_command =>cmd_R42_S146, routeExecute => routes_o(41), clock => clock, reset => reset);
	route_R43 : route_42 port map(routeRequest => routes_i(42), ne17_command => cmd_R43_ne17, track_ne17 => state_ne17, ne59_command => cmd_R43_ne59, track_ne59 => state_ne59, s69W03_command => cmd_R43_69W03, s69W03_state => state_69W03, Sw06_command => cmd_R43_Sw06, Sw06_state => state_Sw06, S83_state => state_S83, S83_command => cmd_R43_S83, C109_state => state_C109, C109_command =>cmd_R43_C109, routeExecute => routes_o(42), clock => clock, reset => reset);
	route_R44 : route_43 port map(routeRequest => routes_i(43), ne11_command => cmd_R44_ne11, track_ne11 => state_ne11, ne59_command => cmd_R44_ne59, track_ne59 => state_ne59, ne95_command => cmd_R44_ne95, track_ne95 => state_ne95, ne52_command => cmd_R44_ne52, track_ne52 => state_ne52, Lc01_command => cmd_R44_Lc01, Lc01_state => state_Lc01, s69W03_command => cmd_R44_69W03, s69W03_state => state_69W03, s69W04_command => cmd_R44_69W04, s69W04_state => state_69W04, S86_state => state_S86, S86_command => cmd_R44_S86, X51_state => state_X51, X51_command =>cmd_R44_X51, routeExecute => routes_o(43), clock => clock, reset => reset);
	route_R45 : route_44 port map(routeRequest => routes_i(44), ne14_command => cmd_R45_ne14, track_ne14 => state_ne14, ne52_command => cmd_R45_ne52, track_ne52 => state_ne52, s69W04_command => cmd_R45_69W04, s69W04_state => state_69W04, S86_state => state_S86, S86_command => cmd_R45_S86, T07_state => state_T07, T07_command =>cmd_R45_T07, routeExecute => routes_o(44), clock => clock, reset => reset);
	route_R46 : route_45 port map(routeRequest => routes_i(45), ne23_command => cmd_R46_ne23, track_ne23 => state_ne23, ne64_command => cmd_R46_ne64, track_ne64 => state_ne64, ne67_command => cmd_R46_ne67, track_ne67 => state_ne67, ne103_command => cmd_R46_ne103, track_ne103 => state_ne103, B89_state => state_B89, B89_command => cmd_R46_B89, P64_state => state_P64, P64_command =>cmd_R46_P64, routeExecute => routes_o(45), clock => clock, reset => reset);
	route_R47 : route_46 port map(routeRequest => routes_i(46), ne23_command => cmd_R47_ne23, track_ne23 => state_ne23, ne64_command => cmd_R47_ne64, track_ne64 => state_ne64, s70W01_command => cmd_R47_70W01, s70W01_state => state_70W01, s70W02_command => cmd_R47_70W02, s70W02_state => state_70W02, S90_state => state_S90, S90_command => cmd_R47_S90, P60_state => state_P60, P60_command =>cmd_R47_P60, routeExecute => routes_o(46), clock => clock, reset => reset);
	route_R48 : route_47 port map(routeRequest => routes_i(47), ne24_command => cmd_R48_ne24, track_ne24 => state_ne24, ne64_command => cmd_R48_ne64, track_ne64 => state_ne64, s70W01_command => cmd_R48_70W01, s70W01_state => state_70W01, s70W02_command => cmd_R48_70W02, s70W02_state => state_70W02, S90_state => state_S90, S90_command => cmd_R48_S90, B92_state => state_B92, B92_command =>cmd_R48_B92, routeExecute => routes_o(47), clock => clock, reset => reset);
	route_R49 : route_48 port map(routeRequest => routes_i(48), ne24_command => cmd_R49_ne24, track_ne24 => state_ne24, ne26_command => cmd_R49_ne26, track_ne26 => state_ne26, s70W02_command => cmd_R49_70W02, s70W02_state => state_70W02, B92_state => state_B92, B92_command => cmd_R49_B92, L27_state => state_L27, L27_command =>cmd_R49_L27, routeExecute => routes_o(48), clock => clock, reset => reset);
	route_R50 : route_49 port map(routeRequest => routes_i(49), ne23_command => cmd_R50_ne23, track_ne23 => state_ne23, ne26_command => cmd_R50_ne26, track_ne26 => state_ne26, s70W02_command => cmd_R50_70W02, s70W02_state => state_70W02, S93_state => state_S93, S93_command => cmd_R50_S93, B89_state => state_B89, B89_command =>cmd_R50_B89, routeExecute => routes_o(49), clock => clock, reset => reset);
	route_R51 : route_50 port map(routeRequest => routes_i(50), ne24_command => cmd_R51_ne24, track_ne24 => state_ne24, ne26_command => cmd_R51_ne26, track_ne26 => state_ne26, s70W02_command => cmd_R51_70W02, s70W02_state => state_70W02, S93_state => state_S93, S93_command => cmd_R51_S93, P63_state => state_P63, P63_command =>cmd_R51_P63, routeExecute => routes_o(50), clock => clock, reset => reset);
	route_R52 : route_51 port map(routeRequest => routes_i(51), ne30_command => cmd_R52_ne30, track_ne30 => state_ne30, ne83_command => cmd_R52_ne83, track_ne83 => state_ne83, Sw08_command => cmd_R52_Sw08, Sw08_state => state_Sw08, Sw12_command => cmd_R52_Sw12, Sw12_state => state_Sw12, C95_state => state_C95, C95_command => cmd_R52_C95, S122_state => state_S122, S122_command =>cmd_R52_S122, routeExecute => routes_o(51), clock => clock, reset => reset);
	route_R53 : route_52 port map(routeRequest => routes_i(52), ne29_command => cmd_R53_ne29, track_ne29 => state_ne29, ne30_command => cmd_R53_ne30, track_ne30 => state_ne30, Sw08_command => cmd_R53_Sw08, Sw08_state => state_Sw08, Sw12_command => cmd_R53_Sw12, Sw12_state => state_Sw12, B96_state => state_B96, B96_command => cmd_R53_B96, S122_state => state_S122, S122_command =>cmd_R53_S122, routeExecute => routes_o(52), clock => clock, reset => reset);
	route_R54 : route_53 port map(routeRequest => routes_i(53), ne29_command => cmd_R54_ne29, track_ne29 => state_ne29, ne30_command => cmd_R54_ne30, track_ne30 => state_ne30, ne110_command => cmd_R54_ne110, track_ne110 => state_ne110, Sw08_command => cmd_R54_Sw08, Sw08_state => state_Sw08, Sw09_command => cmd_R54_Sw09, Sw09_state => state_Sw09, Sw41_command => cmd_R54_Sw41, Sw41_state => state_Sw41, S97_state => state_S97, S97_command => cmd_R54_S97, C138_state => state_C138, C138_command =>cmd_R54_C138, routeExecute => routes_o(53), clock => clock, reset => reset);
	route_R55 : route_54 port map(routeRequest => routes_i(54), ne30_command => cmd_R55_ne30, track_ne30 => state_ne30, ne83_command => cmd_R55_ne83, track_ne83 => state_ne83, Sw08_command => cmd_R55_Sw08, Sw08_state => state_Sw08, Sw04_command => cmd_R55_Sw04, Sw04_state => state_Sw04, S97_state => state_S97, S97_command => cmd_R55_S97, C114_state => state_C114, C114_command =>cmd_R55_C114, routeExecute => routes_o(54), clock => clock, reset => reset);
	route_R56 : route_55 port map(routeRequest => routes_i(55), ne32_command => cmd_R56_ne32, track_ne32 => state_ne32, ne110_command => cmd_R56_ne110, track_ne110 => state_ne110, Sw09_command => cmd_R56_Sw09, Sw09_state => state_Sw09, Sw41_command => cmd_R56_Sw41, Sw41_state => state_Sw41, C100_state => state_C100, C100_command => cmd_R56_C100, C138_state => state_C138, C138_command =>cmd_R56_C138, routeExecute => routes_o(55), clock => clock, reset => reset);
	route_R57 : route_56 port map(routeRequest => routes_i(56), ne29_command => cmd_R57_ne29, track_ne29 => state_ne29, Sw08_command => cmd_R57_Sw08, Sw08_state => state_Sw08, B101_state => state_B101, B101_command => cmd_R57_B101, B96_state => state_B96, B96_command =>cmd_R57_B96, routeExecute => routes_o(56), clock => clock, reset => reset);
	route_R58 : route_57 port map(routeRequest => routes_i(57), ne32_command => cmd_R58_ne32, track_ne32 => state_ne32, ne110_command => cmd_R58_ne110, track_ne110 => state_ne110, Sw09_command => cmd_R58_Sw09, Sw09_state => state_Sw09, Sw04_command => cmd_R58_Sw04, Sw04_state => state_Sw04, S102_state => state_S102, S102_command => cmd_R58_S102, S115_state => state_S115, S115_command =>cmd_R58_S115, routeExecute => routes_o(57), clock => clock, reset => reset);
	route_R59 : route_58 port map(routeRequest => routes_i(58), ne29_command => cmd_R59_ne29, track_ne29 => state_ne29, ne110_command => cmd_R59_ne110, track_ne110 => state_ne110, Sw09_command => cmd_R59_Sw09, Sw09_state => state_Sw09, S102_state => state_S102, S102_command => cmd_R59_S102, B101_state => state_B101, B101_command =>cmd_R59_B101, routeExecute => routes_o(58), clock => clock, reset => reset);
	route_R60 : route_59 port map(routeRequest => routes_i(59), ne44_command => cmd_R60_ne44, track_ne44 => state_ne44, ne102_command => cmd_R60_ne102, track_ne102 => state_ne102, s71W01_command => cmd_R60_71W01, s71W01_state => state_71W01, C104_state => state_C104, C104_command => cmd_R60_C104, L28_state => state_L28, L28_command =>cmd_R60_L28, routeExecute => routes_o(59), clock => clock, reset => reset);
	route_R61 : route_60 port map(routeRequest => routes_i(60), ne43_command => cmd_R61_ne43, track_ne43 => state_ne43, ne44_command => cmd_R61_ne44, track_ne44 => state_ne44, ne48_command => cmd_R61_ne48, track_ne48 => state_ne48, s71W01_command => cmd_R61_71W01, s71W01_state => state_71W01, s71W02_command => cmd_R61_71W02, s71W02_state => state_71W02, S105_state => state_S105, S105_command => cmd_R61_S105, L29_state => state_L29, L29_command =>cmd_R61_L29, routeExecute => routes_o(60), clock => clock, reset => reset);
	route_R62 : route_61 port map(routeRequest => routes_i(61), ne26_command => cmd_R62_ne26, track_ne26 => state_ne26, ne44_command => cmd_R62_ne44, track_ne44 => state_ne44, ne65_command => cmd_R62_ne65, track_ne65 => state_ne65, ne102_command => cmd_R62_ne102, track_ne102 => state_ne102, s70W02_command => cmd_R62_70W02, s70W02_state => state_70W02, s71W01_command => cmd_R62_71W01, s71W01_state => state_71W01, S105_state => state_S105, S105_command => cmd_R62_S105, S93_state => state_S93, S93_command =>cmd_R62_S93, routeExecute => routes_o(61), clock => clock, reset => reset);
	route_R63 : route_62 port map(routeRequest => routes_i(62), ne17_command => cmd_R63_ne17, track_ne17 => state_ne17, ne78_command => cmd_R63_ne78, track_ne78 => state_ne78, Sw06_command => cmd_R63_Sw06, Sw06_state => state_Sw06, C109_state => state_C109, C109_command => cmd_R63_C109, L33_state => state_L33, L33_command =>cmd_R63_L33, routeExecute => routes_o(62), clock => clock, reset => reset);
	route_R64 : route_63 port map(routeRequest => routes_i(63), ne17_command => cmd_R64_ne17, track_ne17 => state_ne17, ne78_command => cmd_R64_ne78, track_ne78 => state_ne78, s69W03_command => cmd_R64_69W03, s69W03_state => state_69W03, Sw06_command => cmd_R64_Sw06, Sw06_state => state_Sw06, S110_state => state_S110, S110_command => cmd_R64_S110, C82_state => state_C82, C82_command =>cmd_R64_C82, routeExecute => routes_o(63), clock => clock, reset => reset);
	route_R65 : route_64 port map(routeRequest => routes_i(64), ne78_command => cmd_R65_ne78, track_ne78 => state_ne78, ne79_command => cmd_R65_ne79, track_ne79 => state_ne79, ne77_command => cmd_R65_ne77, track_ne77 => state_ne77, Sw06_command => cmd_R65_Sw06, Sw06_state => state_Sw06, Sw07_command => cmd_R65_Sw07, Sw07_state => state_Sw07, S110_state => state_S110, S110_command => cmd_R65_S110, B133_state => state_B133, B133_command =>cmd_R65_B133, routeExecute => routes_o(64), clock => clock, reset => reset);
	route_R66 : route_65 port map(routeRequest => routes_i(65), ne78_command => cmd_R66_ne78, track_ne78 => state_ne78, ne79_command => cmd_R66_ne79, track_ne79 => state_ne79, ne21_command => cmd_R66_ne21, track_ne21 => state_ne21, Sw06_command => cmd_R66_Sw06, Sw06_state => state_Sw06, Sw07_command => cmd_R66_Sw07, Sw07_state => state_Sw07, S110_state => state_S110, S110_command => cmd_R66_S110, P72_state => state_P72, P72_command =>cmd_R66_P72, routeExecute => routes_o(65), clock => clock, reset => reset);
	route_R67 : route_66 port map(routeRequest => routes_i(66), ne32_command => cmd_R67_ne32, track_ne32 => state_ne32, ne83_command => cmd_R67_ne83, track_ne83 => state_ne83, Sw09_command => cmd_R67_Sw09, Sw09_state => state_Sw09, Sw04_command => cmd_R67_Sw04, Sw04_state => state_Sw04, C114_state => state_C114, C114_command => cmd_R67_C114, C100_state => state_C100, C100_command =>cmd_R67_C100, routeExecute => routes_o(66), clock => clock, reset => reset);
	route_R68 : route_67 port map(routeRequest => routes_i(67), ne32_command => cmd_R68_ne32, track_ne32 => state_ne32, ne83_command => cmd_R68_ne83, track_ne83 => state_ne83, Sw08_command => cmd_R68_Sw08, Sw08_state => state_Sw08, Sw04_command => cmd_R68_Sw04, Sw04_state => state_Sw04, S115_state => state_S115, S115_command => cmd_R68_S115, C95_state => state_C95, C95_command =>cmd_R68_C95, routeExecute => routes_o(67), clock => clock, reset => reset);
	route_R69 : route_68 port map(routeRequest => routes_i(68), ne32_command => cmd_R69_ne32, track_ne32 => state_ne32, ne41_command => cmd_R69_ne41, track_ne41 => state_ne41, ne82_command => cmd_R69_ne82, track_ne82 => state_ne82, Sw04_command => cmd_R69_Sw04, Sw04_state => state_Sw04, Sw05_command => cmd_R69_Sw05, Sw05_state => state_Sw05, S115_state => state_S115, S115_command => cmd_R69_S115, P58_state => state_P58, P58_command =>cmd_R69_P58, routeExecute => routes_o(68), clock => clock, reset => reset);
	route_R70 : route_69 port map(routeRequest => routes_i(69), ne32_command => cmd_R70_ne32, track_ne32 => state_ne32, ne82_command => cmd_R70_ne82, track_ne82 => state_ne82, ne84_command => cmd_R70_ne84, track_ne84 => state_ne84, Sw04_command => cmd_R70_Sw04, Sw04_state => state_Sw04, Sw05_command => cmd_R70_Sw05, Sw05_state => state_Sw05, S115_state => state_S115, S115_command => cmd_R70_S115, T13_state => state_T13, T13_command =>cmd_R70_T13, routeExecute => routes_o(69), clock => clock, reset => reset);
	route_R71 : route_70 port map(routeRequest => routes_i(70), ne86_command => cmd_R71_ne86, track_ne86 => state_ne86, ne88_command => cmd_R71_ne88, track_ne88 => state_ne88, Sw11_command => cmd_R71_Sw11, Sw11_state => state_Sw11, C118_state => state_C118, C118_command => cmd_R71_C118, T15_state => state_T15, T15_command =>cmd_R71_T15, routeExecute => routes_o(70), clock => clock, reset => reset);
	route_R72 : route_71 port map(routeRequest => routes_i(71), ne86_command => cmd_R72_ne86, track_ne86 => state_ne86, ne88_command => cmd_R72_ne88, track_ne88 => state_ne88, Sw11_command => cmd_R72_Sw11, Sw11_state => state_Sw11, S119_state => state_S119, S119_command => cmd_R72_S119, T17_state => state_T17, T17_command =>cmd_R72_T17, routeExecute => routes_o(71), clock => clock, reset => reset);
	route_R73 : route_72 port map(routeRequest => routes_i(72), ne30_command => cmd_R73_ne30, track_ne30 => state_ne30, ne86_command => cmd_R73_ne86, track_ne86 => state_ne86, ne87_command => cmd_R73_ne87, track_ne87 => state_ne87, ne91_command => cmd_R73_ne91, track_ne91 => state_ne91, Sw08_command => cmd_R73_Sw08, Sw08_state => state_Sw08, Sw09_command => cmd_R73_Sw09, Sw09_state => state_Sw09, Sw12_command => cmd_R73_Sw12, Sw12_state => state_Sw12, Sw11_command => cmd_R73_Sw11, Sw11_state => state_Sw11, Sw13_command => cmd_R73_Sw13, Sw13_state => state_Sw13, S119_state => state_S119, S119_command => cmd_R73_S119, S97_state => state_S97, S97_command =>cmd_R73_S97, routeExecute => routes_o(72), clock => clock, reset => reset);
	route_R74 : route_73 port map(routeRequest => routes_i(73), ne30_command => cmd_R74_ne30, track_ne30 => state_ne30, ne89_command => cmd_R74_ne89, track_ne89 => state_ne89, Sw12_command => cmd_R74_Sw12, Sw12_state => state_Sw12, S122_state => state_S122, S122_command => cmd_R74_S122, T19_state => state_T19, T19_command =>cmd_R74_T19, routeExecute => routes_o(73), clock => clock, reset => reset);
	route_R75 : route_74 port map(routeRequest => routes_i(74), ne30_command => cmd_R75_ne30, track_ne30 => state_ne30, ne86_command => cmd_R75_ne86, track_ne86 => state_ne86, ne87_command => cmd_R75_ne87, track_ne87 => state_ne87, ne91_command => cmd_R75_ne91, track_ne91 => state_ne91, Sw12_command => cmd_R75_Sw12, Sw12_state => state_Sw12, Sw11_command => cmd_R75_Sw11, Sw11_state => state_Sw11, Sw13_command => cmd_R75_Sw13, Sw13_state => state_Sw13, S122_state => state_S122, S122_command => cmd_R75_S122, T15_state => state_T15, T15_command =>cmd_R75_T15, routeExecute => routes_o(74), clock => clock, reset => reset);
	route_R76 : route_75 port map(routeRequest => routes_i(75), ne30_command => cmd_R76_ne30, track_ne30 => state_ne30, ne90_command => cmd_R76_ne90, track_ne90 => state_ne90, ne91_command => cmd_R76_ne91, track_ne91 => state_ne91, Sw12_command => cmd_R76_Sw12, Sw12_state => state_Sw12, Sw13_command => cmd_R76_Sw13, Sw13_state => state_Sw13, S122_state => state_S122, S122_command => cmd_R76_S122, T21_state => state_T21, T21_command =>cmd_R76_T21, routeExecute => routes_o(75), clock => clock, reset => reset);
	route_R77 : route_76 port map(routeRequest => routes_i(76), ne32_command => cmd_R77_ne32, track_ne32 => state_ne32, ne41_command => cmd_R77_ne41, track_ne41 => state_ne41, ne82_command => cmd_R77_ne82, track_ne82 => state_ne82, Sw09_command => cmd_R77_Sw09, Sw09_state => state_Sw09, Sw04_command => cmd_R77_Sw04, Sw04_state => state_Sw04, Sw05_command => cmd_R77_Sw05, Sw05_state => state_Sw05, B130_state => state_B130, B130_command => cmd_R77_B130, C100_state => state_C100, C100_command =>cmd_R77_C100, routeExecute => routes_o(76), clock => clock, reset => reset);
	route_R78 : route_77 port map(routeRequest => routes_i(77), ne41_command => cmd_R78_ne41, track_ne41 => state_ne41, ne44_command => cmd_R78_ne44, track_ne44 => state_ne44, ne100_command => cmd_R78_ne100, track_ne100 => state_ne100, ne101_command => cmd_R78_ne101, track_ne101 => state_ne101, ne85_command => cmd_R78_ne85, track_ne85 => state_ne85, s71W01_command => cmd_R78_71W01, s71W01_state => state_71W01, s71W02_command => cmd_R78_71W02, s71W02_state => state_71W02, Sw41_command => cmd_R78_Sw41, Sw41_state => state_Sw41, Sw05_command => cmd_R78_Sw05, Sw05_state => state_Sw05, B130_state => state_B130, B130_command => cmd_R78_B130, S105_state => state_S105, S105_command =>cmd_R78_S105, routeExecute => routes_o(77), clock => clock, reset => reset);
	route_R79 : route_78 port map(routeRequest => routes_i(78), ne41_command => cmd_R79_ne41, track_ne41 => state_ne41, ne85_command => cmd_R79_ne85, track_ne85 => state_ne85, Sw05_command => cmd_R79_Sw05, Sw05_state => state_Sw05, S131_state => state_S131, S131_command => cmd_R79_S131, P58_state => state_P58, P58_command =>cmd_R79_P58, routeExecute => routes_o(78), clock => clock, reset => reset);
	route_R80 : route_79 port map(routeRequest => routes_i(79), ne84_command => cmd_R80_ne84, track_ne84 => state_ne84, ne85_command => cmd_R80_ne85, track_ne85 => state_ne85, Sw05_command => cmd_R80_Sw05, Sw05_state => state_Sw05, S131_state => state_S131, S131_command => cmd_R80_S131, T13_state => state_T13, T13_command =>cmd_R80_T13, routeExecute => routes_o(79), clock => clock, reset => reset);
	route_R81 : route_80 port map(routeRequest => routes_i(80), ne77_command => cmd_R81_ne77, track_ne77 => state_ne77, ne52_command => cmd_R81_ne52, track_ne52 => state_ne52, s69W03_command => cmd_R81_69W03, s69W03_state => state_69W03, s69W04_command => cmd_R81_69W04, s69W04_state => state_69W04, Sw03_command => cmd_R81_Sw03, Sw03_state => state_Sw03, B133_state => state_B133, B133_command => cmd_R81_B133, S86_state => state_S86, S86_command =>cmd_R81_S86, routeExecute => routes_o(80), clock => clock, reset => reset);
	route_R82 : route_81 port map(routeRequest => routes_i(81), ne94_command => cmd_R82_ne94, track_ne94 => state_ne94, ne77_command => cmd_R82_ne77, track_ne77 => state_ne77, Sw07_command => cmd_R82_Sw07, Sw07_state => state_Sw07, S135_state => state_S135, S135_command => cmd_R82_S135, B133_state => state_B133, B133_command =>cmd_R82_B133, routeExecute => routes_o(81), clock => clock, reset => reset);
	route_R83 : route_82 port map(routeRequest => routes_i(82), ne94_command => cmd_R83_ne94, track_ne94 => state_ne94, ne21_command => cmd_R83_ne21, track_ne21 => state_ne21, Sw07_command => cmd_R83_Sw07, Sw07_state => state_Sw07, S135_state => state_S135, S135_command => cmd_R83_S135, P72_state => state_P72, P72_command =>cmd_R83_P72, routeExecute => routes_o(82), clock => clock, reset => reset);
	route_R84 : route_83 port map(routeRequest => routes_i(83), ne44_command => cmd_R84_ne44, track_ne44 => state_ne44, ne100_command => cmd_R84_ne100, track_ne100 => state_ne100, ne101_command => cmd_R84_ne101, track_ne101 => state_ne101, ne110_command => cmd_R84_ne110, track_ne110 => state_ne110, s71W01_command => cmd_R84_71W01, s71W01_state => state_71W01, s71W02_command => cmd_R84_71W02, s71W02_state => state_71W02, Sw41_command => cmd_R84_Sw41, Sw41_state => state_Sw41, C138_state => state_C138, C138_command => cmd_R84_C138, S105_state => state_S105, S105_command =>cmd_R84_S105, routeExecute => routes_o(83), clock => clock, reset => reset);
	route_R85 : route_84 port map(routeRequest => routes_i(84), ne100_command => cmd_R85_ne100, track_ne100 => state_ne100, ne110_command => cmd_R85_ne110, track_ne110 => state_ne110, Sw09_command => cmd_R85_Sw09, Sw09_state => state_Sw09, Sw41_command => cmd_R85_Sw41, Sw41_state => state_Sw41, S139_state => state_S139, S139_command => cmd_R85_S139, S102_state => state_S102, S102_command =>cmd_R85_S102, routeExecute => routes_o(84), clock => clock, reset => reset);
	route_R86 : route_85 port map(routeRequest => routes_i(85), ne100_command => cmd_R86_ne100, track_ne100 => state_ne100, ne85_command => cmd_R86_ne85, track_ne85 => state_ne85, Sw41_command => cmd_R86_Sw41, Sw41_state => state_Sw41, S139_state => state_S139, S139_command => cmd_R86_S139, S131_state => state_S131, S131_command =>cmd_R86_S131, routeExecute => routes_o(85), clock => clock, reset => reset);
	route_R87 : route_86 port map(routeRequest => routes_i(86), ne70_command => cmd_R87_ne70, track_ne70 => state_ne70, ne104_command => cmd_R87_ne104, track_ne104 => state_ne104, B143_state => state_B143, B143_command => cmd_R87_B143, L32_state => state_L32, L32_command =>cmd_R87_L32, routeExecute => routes_o(86), clock => clock, reset => reset);
	route_R88 : route_87 port map(routeRequest => routes_i(87), ne104_command => cmd_R88_ne104, track_ne104 => state_ne104, ne21_command => cmd_R88_ne21, track_ne21 => state_ne21, Sw03_command => cmd_R88_Sw03, Sw03_state => state_Sw03, S144_state => state_S144, S144_command => cmd_R88_S144, B143_state => state_B143, B143_command =>cmd_R88_B143, routeExecute => routes_o(87), clock => clock, reset => reset);
	route_R89 : route_88 port map(routeRequest => routes_i(88), ne78_command => cmd_R89_ne78, track_ne78 => state_ne78, ne79_command => cmd_R89_ne79, track_ne79 => state_ne79, ne77_command => cmd_R89_ne77, track_ne77 => state_ne77, Sw06_command => cmd_R89_Sw06, Sw06_state => state_Sw06, Sw07_command => cmd_R89_Sw07, Sw07_state => state_Sw07, B145_state => state_B145, B145_command => cmd_R89_B145, L33_state => state_L33, L33_command =>cmd_R89_L33, routeExecute => routes_o(88), clock => clock, reset => reset);
	route_R90 : route_89 port map(routeRequest => routes_i(89), ne94_command => cmd_R90_ne94, track_ne94 => state_ne94, ne97_command => cmd_R90_ne97, track_ne97 => state_ne97, ne99_command => cmd_R90_ne99, track_ne99 => state_ne99, ne77_command => cmd_R90_ne77, track_ne77 => state_ne77, Sw07_command => cmd_R90_Sw07, Sw07_state => state_Sw07, B145_state => state_B145, B145_command => cmd_R90_B145, P69_state => state_P69, P69_command =>cmd_R90_P69, routeExecute => routes_o(89), clock => clock, reset => reset);
	route_R91 : route_90 port map(routeRequest => routes_i(90), ne77_command => cmd_R91_ne77, track_ne77 => state_ne77, ne52_command => cmd_R91_ne52, track_ne52 => state_ne52, Sw06_command => cmd_R91_Sw06, Sw06_state => state_Sw06, Sw03_command => cmd_R91_Sw03, Sw03_state => state_Sw03, S146_state => state_S146, S146_command => cmd_R91_S146, B145_state => state_B145, B145_command =>cmd_R91_B145, routeExecute => routes_o(90), clock => clock, reset => reset);
	processed <= processing;
	tracks_o(0) <= state_ne1;
	tracks_o(1) <= state_ne4;
	tracks_o(2) <= state_ne7;
	tracks_o(3) <= state_ne9;
	tracks_o(4) <= state_ne11;
	tracks_o(5) <= state_ne14;
	tracks_o(6) <= state_ne17;
	tracks_o(7) <= state_ne23;
	tracks_o(8) <= state_ne24;
	tracks_o(9) <= state_ne26;
	tracks_o(10) <= state_ne29;
	tracks_o(11) <= state_ne30;
	tracks_o(12) <= state_ne32;
	tracks_o(13) <= state_ne41;
	tracks_o(14) <= state_ne43;
	tracks_o(15) <= state_ne44;
	tracks_o(16) <= state_ne47;
	tracks_o(17) <= state_ne48;
	tracks_o(18) <= state_ne59;
	tracks_o(19) <= state_ne64;
	tracks_o(20) <= state_ne65;
	tracks_o(21) <= state_ne67;
	tracks_o(22) <= state_ne70;
	tracks_o(23) <= state_ne78;
	tracks_o(24) <= state_ne79;
	tracks_o(25) <= state_ne82;
	tracks_o(26) <= state_ne83;
	tracks_o(27) <= state_ne84;
	tracks_o(28) <= state_ne86;
	tracks_o(29) <= state_ne87;
	tracks_o(30) <= state_ne88;
	tracks_o(31) <= state_ne89;
	tracks_o(32) <= state_ne90;
	tracks_o(33) <= state_ne91;
	tracks_o(34) <= state_ne93;
	tracks_o(35) <= state_ne94;
	tracks_o(36) <= state_ne95;
	tracks_o(37) <= state_ne96;
	tracks_o(38) <= state_ne97;
	tracks_o(39) <= state_ne98;
	tracks_o(40) <= state_ne99;
	tracks_o(41) <= state_ne100;
	tracks_o(42) <= state_ne101;
	tracks_o(43) <= state_ne102;
	tracks_o(44) <= state_ne103;
	tracks_o(45) <= state_ne105;
	tracks_o(46) <= state_ne106;
	tracks_o(47) <= state_ne85;
	tracks_o(48) <= state_ne77;
	tracks_o(49) <= state_ne104;
	tracks_o(50) <= state_ne52;
	tracks_o(51) <= state_ne21;
	tracks_o(52) <= state_ne110;
end Behavioral;