--  splitter.vhdl : Automatically generated using ACG
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
--Declare the package
use work.my_package.all;
	entity splitter is
		generic(
			N : natural := 329;
			N_SIGNALS : natural := 82;
			N_LEVELCROSSINGS : natural := 1;
			N_SINGLESWITCHES : natural := 15;
			N_DOUBLEWITCHES : natural := 2;
			N_SCRISSORCROSSINGS : natural := 1;
			N_ROUTES : natural := 91;
			N_TRACKCIRCUITS : natural := 53
		);
		port(
			clock : in std_logic;
			packet :  in std_logic_vector(N-1 downto 0);
			processing :  in std_logic;
			processed :  out std_logic;
			ocupation :  out std_logic_vector(N_TRACKCIRCUITS-1 downto 0);
			signals :  out signals_type;
			routes : out std_logic_vector(N_ROUTES-1 downto 0);
			levelCrossings : out std_logic;
			singleSwitches : out std_logic_vector(N_SINGLESWITCHES-1 downto 0);
			scissorSwitches : out std_logic;
			doubleSwitches : out dSwitches_type;
			reset : in std_logic
		);
	end entity splitter;
architecture Behavioral of splitter is
	Signal tc_s : std_logic_vector(53-1 downto 0);
	Signal sig_s_i,sig_s_o : signals_type;
	Signal rt_s_i,rt_s_o : std_logic_vector(91-1 downto 0);
	Signal lc_s_i,lc_s_o : std_logic;
	Signal ssw_s_i,ssw_s_o : std_logic_vector(15-1 downto 0);
	Signal sc_s_i,sc_s_o : std_logic;
	Signal dsw_s_i,dsw_s_o : dSwitches_type;
begin
	process(clock,reset)
	begin
		if (clock = '1' and clock'Event) then
			if (reset = '1') then
				ocupation <= "00000000000000000000000000000000000000000000000000000";
				signals.lsb <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000";
				signals.msb <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000";
				routes <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
				levelCrossings <= '0';
				singleSwitches <= "000000000000000";
				scissorSwitches <= '0';
				doubleSwitches.lsb <= "00";
				doubleSwitches.msb <= "00";
				processed <= '0';
			else
				processed <= processing;
				if processing = '1' then
					ocupation(0) <= packet(328);
					ocupation(1) <= packet(327);
					ocupation(2) <= packet(326);
					ocupation(3) <= packet(325);
					ocupation(4) <= packet(324);
					ocupation(5) <= packet(323);
					ocupation(6) <= packet(322);
					ocupation(7) <= packet(321);
					ocupation(8) <= packet(320);
					ocupation(9) <= packet(319);
					ocupation(10) <= packet(318);
					ocupation(11) <= packet(317);
					ocupation(12) <= packet(316);
					ocupation(13) <= packet(315);
					ocupation(14) <= packet(314);
					ocupation(15) <= packet(313);
					ocupation(16) <= packet(312);
					ocupation(17) <= packet(311);
					ocupation(18) <= packet(310);
					ocupation(19) <= packet(309);
					ocupation(20) <= packet(308);
					ocupation(21) <= packet(307);
					ocupation(22) <= packet(306);
					ocupation(23) <= packet(305);
					ocupation(24) <= packet(304);
					ocupation(25) <= packet(303);
					ocupation(26) <= packet(302);
					ocupation(27) <= packet(301);
					ocupation(28) <= packet(300);
					ocupation(29) <= packet(299);
					ocupation(30) <= packet(298);
					ocupation(31) <= packet(297);
					ocupation(32) <= packet(296);
					ocupation(33) <= packet(295);
					ocupation(34) <= packet(294);
					ocupation(35) <= packet(293);
					ocupation(36) <= packet(292);
					ocupation(37) <= packet(291);
					ocupation(38) <= packet(290);
					ocupation(39) <= packet(289);
					ocupation(40) <= packet(288);
					ocupation(41) <= packet(287);
					ocupation(42) <= packet(286);
					ocupation(43) <= packet(285);
					ocupation(44) <= packet(284);
					ocupation(45) <= packet(283);
					ocupation(46) <= packet(282);
					ocupation(47) <= packet(281);
					ocupation(48) <= packet(280);
					ocupation(49) <= packet(279);
					ocupation(50) <= packet(278);
					ocupation(51) <= packet(277);
					ocupation(52) <= packet(276);
					routes(0) <= packet(275);
					routes(1) <= packet(274);
					routes(2) <= packet(273);
					routes(3) <= packet(272);
					routes(4) <= packet(271);
					routes(5) <= packet(270);
					routes(6) <= packet(269);
					routes(7) <= packet(268);
					routes(8) <= packet(267);
					routes(9) <= packet(266);
					routes(10) <= packet(265);
					routes(11) <= packet(264);
					routes(12) <= packet(263);
					routes(13) <= packet(262);
					routes(14) <= packet(261);
					routes(15) <= packet(260);
					routes(16) <= packet(259);
					routes(17) <= packet(258);
					routes(18) <= packet(257);
					routes(19) <= packet(256);
					routes(20) <= packet(255);
					routes(21) <= packet(254);
					routes(22) <= packet(253);
					routes(23) <= packet(252);
					routes(24) <= packet(251);
					routes(25) <= packet(250);
					routes(26) <= packet(249);
					routes(27) <= packet(248);
					routes(28) <= packet(247);
					routes(29) <= packet(246);
					routes(30) <= packet(245);
					routes(31) <= packet(244);
					routes(32) <= packet(243);
					routes(33) <= packet(242);
					routes(34) <= packet(241);
					routes(35) <= packet(240);
					routes(36) <= packet(239);
					routes(37) <= packet(238);
					routes(38) <= packet(237);
					routes(39) <= packet(236);
					routes(40) <= packet(235);
					routes(41) <= packet(234);
					routes(42) <= packet(233);
					routes(43) <= packet(232);
					routes(44) <= packet(231);
					routes(45) <= packet(230);
					routes(46) <= packet(229);
					routes(47) <= packet(228);
					routes(48) <= packet(227);
					routes(49) <= packet(226);
					routes(50) <= packet(225);
					routes(51) <= packet(224);
					routes(52) <= packet(223);
					routes(53) <= packet(222);
					routes(54) <= packet(221);
					routes(55) <= packet(220);
					routes(56) <= packet(219);
					routes(57) <= packet(218);
					routes(58) <= packet(217);
					routes(59) <= packet(216);
					routes(60) <= packet(215);
					routes(61) <= packet(214);
					routes(62) <= packet(213);
					routes(63) <= packet(212);
					routes(64) <= packet(211);
					routes(65) <= packet(210);
					routes(66) <= packet(209);
					routes(67) <= packet(208);
					routes(68) <= packet(207);
					routes(69) <= packet(206);
					routes(70) <= packet(205);
					routes(71) <= packet(204);
					routes(72) <= packet(203);
					routes(73) <= packet(202);
					routes(74) <= packet(201);
					routes(75) <= packet(200);
					routes(76) <= packet(199);
					routes(77) <= packet(198);
					routes(78) <= packet(197);
					routes(79) <= packet(196);
					routes(80) <= packet(195);
					routes(81) <= packet(194);
					routes(82) <= packet(193);
					routes(83) <= packet(192);
					routes(84) <= packet(191);
					routes(85) <= packet(190);
					routes(86) <= packet(189);
					routes(87) <= packet(188);
					routes(88) <= packet(187);
					routes(89) <= packet(186);
					routes(90) <= packet(185);
					signals.msb(0) <= packet(184);
					signals.lsb(0) <= packet(183);
					signals.msb(1) <= packet(182);
					signals.lsb(1) <= packet(181);
					signals.msb(2) <= packet(180);
					signals.lsb(2) <= packet(179);
					signals.msb(3) <= packet(178);
					signals.lsb(3) <= packet(177);
					signals.msb(4) <= packet(176);
					signals.lsb(4) <= packet(175);
					signals.msb(5) <= packet(174);
					signals.lsb(5) <= packet(173);
					signals.msb(6) <= packet(172);
					signals.lsb(6) <= packet(171);
					signals.msb(7) <= packet(170);
					signals.lsb(7) <= packet(169);
					signals.msb(8) <= packet(168);
					signals.lsb(8) <= packet(167);
					signals.msb(9) <= packet(166);
					signals.lsb(9) <= packet(165);
					signals.msb(10) <= packet(164);
					signals.lsb(10) <= packet(163);
					signals.msb(11) <= packet(162);
					signals.lsb(11) <= packet(161);
					signals.msb(12) <= packet(160);
					signals.lsb(12) <= packet(159);
					signals.msb(13) <= packet(158);
					signals.lsb(13) <= packet(157);
					signals.msb(14) <= packet(156);
					signals.lsb(14) <= packet(155);
					signals.msb(15) <= packet(154);
					signals.lsb(15) <= packet(153);
					signals.msb(16) <= packet(152);
					signals.lsb(16) <= packet(151);
					signals.msb(17) <= packet(150);
					signals.lsb(17) <= packet(149);
					signals.msb(18) <= packet(148);
					signals.lsb(18) <= packet(147);
					signals.msb(19) <= packet(146);
					signals.lsb(19) <= packet(145);
					signals.msb(20) <= packet(144);
					signals.lsb(20) <= packet(143);
					signals.msb(21) <= packet(142);
					signals.lsb(21) <= packet(141);
					signals.msb(22) <= packet(140);
					signals.lsb(22) <= packet(139);
					signals.msb(23) <= packet(138);
					signals.lsb(23) <= packet(137);
					signals.msb(24) <= packet(136);
					signals.lsb(24) <= packet(135);
					signals.msb(25) <= packet(134);
					signals.lsb(25) <= packet(133);
					signals.msb(26) <= packet(132);
					signals.lsb(26) <= packet(131);
					signals.msb(27) <= packet(130);
					signals.lsb(27) <= packet(129);
					signals.msb(28) <= packet(128);
					signals.lsb(28) <= packet(127);
					signals.msb(29) <= packet(126);
					signals.lsb(29) <= packet(125);
					signals.msb(30) <= packet(124);
					signals.lsb(30) <= packet(123);
					signals.msb(31) <= packet(122);
					signals.lsb(31) <= packet(121);
					signals.msb(32) <= packet(120);
					signals.lsb(32) <= packet(119);
					signals.msb(33) <= packet(118);
					signals.lsb(33) <= packet(117);
					signals.msb(34) <= packet(116);
					signals.lsb(34) <= packet(115);
					signals.msb(35) <= packet(114);
					signals.lsb(35) <= packet(113);
					signals.msb(36) <= packet(112);
					signals.lsb(36) <= packet(111);
					signals.msb(37) <= packet(110);
					signals.lsb(37) <= packet(109);
					signals.msb(38) <= packet(108);
					signals.lsb(38) <= packet(107);
					signals.msb(39) <= packet(106);
					signals.lsb(39) <= packet(105);
					signals.msb(40) <= packet(104);
					signals.lsb(40) <= packet(103);
					signals.msb(41) <= packet(102);
					signals.lsb(41) <= packet(101);
					signals.msb(42) <= packet(100);
					signals.lsb(42) <= packet(99);
					signals.msb(43) <= packet(98);
					signals.lsb(43) <= packet(97);
					signals.msb(44) <= packet(96);
					signals.lsb(44) <= packet(95);
					signals.msb(45) <= packet(94);
					signals.lsb(45) <= packet(93);
					signals.msb(46) <= packet(92);
					signals.lsb(46) <= packet(91);
					signals.msb(47) <= packet(90);
					signals.lsb(47) <= packet(89);
					signals.msb(48) <= packet(88);
					signals.lsb(48) <= packet(87);
					signals.msb(49) <= packet(86);
					signals.lsb(49) <= packet(85);
					signals.msb(50) <= packet(84);
					signals.lsb(50) <= packet(83);
					signals.msb(51) <= packet(82);
					signals.lsb(51) <= packet(81);
					signals.msb(52) <= packet(80);
					signals.lsb(52) <= packet(79);
					signals.msb(53) <= packet(78);
					signals.lsb(53) <= packet(77);
					signals.msb(54) <= packet(76);
					signals.lsb(54) <= packet(75);
					signals.msb(55) <= packet(74);
					signals.lsb(55) <= packet(73);
					signals.msb(56) <= packet(72);
					signals.lsb(56) <= packet(71);
					signals.msb(57) <= packet(70);
					signals.lsb(57) <= packet(69);
					signals.msb(58) <= packet(68);
					signals.lsb(58) <= packet(67);
					signals.msb(59) <= packet(66);
					signals.lsb(59) <= packet(65);
					signals.msb(60) <= packet(64);
					signals.lsb(60) <= packet(63);
					signals.msb(61) <= packet(62);
					signals.lsb(61) <= packet(61);
					signals.msb(62) <= packet(60);
					signals.lsb(62) <= packet(59);
					signals.msb(63) <= packet(58);
					signals.lsb(63) <= packet(57);
					signals.msb(64) <= packet(56);
					signals.lsb(64) <= packet(55);
					signals.msb(65) <= packet(54);
					signals.lsb(65) <= packet(53);
					signals.msb(66) <= packet(52);
					signals.lsb(66) <= packet(51);
					signals.msb(67) <= packet(50);
					signals.lsb(67) <= packet(49);
					signals.msb(68) <= packet(48);
					signals.lsb(68) <= packet(47);
					signals.msb(69) <= packet(46);
					signals.lsb(69) <= packet(45);
					signals.msb(70) <= packet(44);
					signals.lsb(70) <= packet(43);
					signals.msb(71) <= packet(42);
					signals.lsb(71) <= packet(41);
					signals.msb(72) <= packet(40);
					signals.lsb(72) <= packet(39);
					signals.msb(73) <= packet(38);
					signals.lsb(73) <= packet(37);
					signals.msb(74) <= packet(36);
					signals.lsb(74) <= packet(35);
					signals.msb(75) <= packet(34);
					signals.lsb(75) <= packet(33);
					signals.msb(76) <= packet(32);
					signals.lsb(76) <= packet(31);
					signals.msb(77) <= packet(30);
					signals.lsb(77) <= packet(29);
					signals.msb(78) <= packet(28);
					signals.lsb(78) <= packet(27);
					signals.msb(79) <= packet(26);
					signals.lsb(79) <= packet(25);
					signals.msb(80) <= packet(24);
					signals.lsb(80) <= packet(23);
					signals.msb(81) <= packet(22);
					signals.lsb(81) <= packet(21);
					levelCrossings <= packet(20);
					singleSwitches(0) <= packet(19);
					singleSwitches(1) <= packet(18);
					singleSwitches(2) <= packet(17);
					singleSwitches(3) <= packet(16);
					singleSwitches(4) <= packet(15);
					singleSwitches(5) <= packet(14);
					singleSwitches(6) <= packet(13);
					singleSwitches(7) <= packet(12);
					singleSwitches(8) <= packet(11);
					singleSwitches(9) <= packet(10);
					singleSwitches(10) <= packet(9);
					singleSwitches(11) <= packet(8);
					singleSwitches(12) <= packet(7);
					singleSwitches(13) <= packet(6);
					singleSwitches(14) <= packet(5);
					doubleSwitches.msb(0) <= packet(4);
					doubleSwitches.lsb(0) <= packet(3);
					doubleSwitches.msb(1) <= packet(2);
					doubleSwitches.lsb(1) <= packet(1);
					scissorCrossings <= packet(-1);
				end if;
			end if;
		end if;
	end process;
end Behavioral;